"Vi har nu 4 månader gamla möss som är icke-diabetiker som brukade vara diabetiker", tillade han.
Dr Ehud Ur, professor i medicin vid Dalhousie University i Halifax, Nova Scotia och ordförande för den kliniska och vetenskapliga avdelningen av Canadian Diabetes Association varnade för att forskningen fortfarande är i sin linda.
Liksom vissa andra experter är han skeptisk till om diabetes kan botas och noterar att dessa fynd inte har någon relevans för personer som redan har typ 1-diabetes.
I måndags meddelade Sara Danius, ständig sekreterare i Svenska Akademiens Nobelkommitté för litteratur, i ett radioprogram i Sveriges Radio att kommittén, som inte kunde nå Bob Dylan direkt om att vinna Nobelpriset i litteratur 2016, hade gett upp sina försök att nå honom.
Danius svarade: "Just nu gör vi ingenting. Jag har ringt och skickat e-post till hans närmaste samarbetspartner och fått mycket vänliga svar. För tillfället räcker det verkligen."
Tidigare har Rings VD, Jamie Siminoff, påpekat att företaget startade när hans dörrklocka inte hördes från hans butik i hans garage.
Han byggde en WiFi-dörrklocka, sa han.
Siminoff sa att försäljningen ökade efter hans framträdande 2013 i ett Shark Tank-avsnitt där showpanelen avböjde att finansiera startupen.
I slutet av 2017 dök Siminoff upp på shopping-tv-kanalen QVC.
Ring gjorde också upp med det konkurrerande säkerhetsföretaget ADT Corporation.
Även om ett experimentellt vaccin verkar kunna minska dödligheten i ebola, har hittills inga läkemedel tydligt visat sig vara lämpliga för att behandla befintliga infektioner.
En antikroppscocktail, ZMapp, visade sig till en början lovande inom området, men formella studier visade att den hade mindre nytta än vad som eftersträvades för att förhindra dödsfall.
I PALM-studien fungerade ZMapp som en kontroll, vilket innebär att forskarna använde den som en baslinje och jämförde de tre andra behandlingarna med den.
USA Gymnastics stöder USA:s olympiska kommittés brev och accepterar det absoluta behovet av den olympiska familjen för att främja en säker miljö för alla våra idrottare.
Vi håller med USOC:s uttalande om att våra idrottares och klubbars intressen, och deras sport, kan tjänas bättre genom att gå vidare med meningsfulla förändringar inom vår organisation, snarare än avcertifiering.
USA Gymnastics stöder en oberoende utredning som kan belysa hur övergrepp av den omfattning som så modigt beskrivits av de överlevande från Larry Nassar kunde ha gått oupptäckt under så lång tid och omfattar alla nödvändiga och lämpliga förändringar.
USA Gymnastics och USOC har samma mål - att göra gymnastiksporten och andra så säkra som möjligt för idrottare att följa sina drömmar i en säker, positiv och bemyndigad miljö.
Under hela 1960-talet arbetade Brzezinski för John F. Kennedy som hans rådgivare och sedan för Lyndon B. Johnsons administration.
Under valet 1976 var han rådgivare till Carter i utrikespolitik och tjänstgjorde sedan som nationell säkerhetsrådgivare (NSA) från 1977 till 1981, där han efterträdde Henry Kissinger.
Som NSA hjälpte han Carter att diplomatiskt hantera världsfrågor, såsom Camp David-avtalen, 1978; normalisera relationerna mellan USA och Kina i slutet av 1970-talet; den iranska revolutionen, som ledde till gisslankrisen i Iran, 1979; och den sovjetiska invasionen i Afghanistan 1979.
Filmen, med Ryan Gosling och Emma Stone i huvudrollerna, fick nomineringar i alla större kategorier.
Gosling och Stone fick nomineringar för bästa manliga huvudroll respektive skådespelerska.
De övriga nomineringarna inkluderar bästa film, regi, foto, kostymdesign, filmklippning, originalmusik, produktionsdesign, ljudredigering, ljudmixning och originalmanus.
Två låtar från filmen, Audition (The Fools Who Dream) och City of Stars, nominerades för bästa originalsång. Lionsgate-studion fick 26 nomineringar – fler än någon annan studio.
Sent på söndagen meddelade USA:s president Donald Trump i ett uttalande via pressekreteraren att amerikanska trupper kommer att lämna Syrien.
Tillkännagivandet gjordes efter att Trump haft ett telefonsamtal med Turkiets president Recep Tayyip Erdoğan.
Turkiet skulle också ta över bevakningen av tillfångatagna IS-krigare, som europeiska nationer har vägrat att repatriera.
Detta bekräftar inte bara att åtminstone vissa dinosaurier hade fjädrar, en teori som redan är utbredd, utan ger också detaljer som fossil i allmänhet inte kan, såsom färg och tredimensionellt arrangemang.
. Forskare säger att detta djurs fjäderdräkt var kastanjebrun på ovansidan med en blek eller karotenoidfärgad undersida.
Fyndet ger också en inblick i hur fjädrar har utvecklats hos fåglar.
Eftersom dinosauriernas fjädrar inte har ett välutvecklat skaft, en så kallad rachis, men har andra egenskaper hos fjädrar - hullingar och hullingar - drog forskarna slutsatsen att rachis sannolikt var en senare evolutionär utveckling än dessa andra egenskaper.
Fjädrarnas struktur tyder på att de inte användes under flygning utan snarare för temperaturreglering eller uppvisning. Forskarna föreslog att även om detta är svansen på en ung dinosaurie, visar provet vuxen fjäderdräkt och inte en unges dun.
Forskarna föreslog att även om detta är svansen på en ung dinosaurie, visar provet vuxen fjäderdräkt och inte en unges dun.
En bilbomb som detonerade vid polishögkvarteret i Gaziantep, Turkiet i går morse, dödade två poliser och skadade mer än tjugo andra personer.
Guvernörens kontor sade att nitton av de skadade var poliser.
Polisen uppger att de misstänker att en påstådd militant medlem av Daesh (ISIL) är ansvarig för attacken.
De fann att solen fungerade enligt samma grundläggande principer som andra stjärnor: Aktiviteten hos alla stjärnor i systemet visade sig drivas av deras luminositet, deras rotation och inget annat.
Luminositeten och rotationen används tillsammans för att bestämma en stjärnas Rossby-tal, som är relaterat till plasmaflödet.
Ju mindre Rossby-talet är, desto mindre aktiv är stjärnan med avseende på magnetiska omkastningar.
Under sin resa stötte Iwasaki på problem vid många tillfällen.
Han rånades av pirater, attackerades i Tibet av en rabiessmittad hund, flydde från äktenskap i Nepal och arresterades i Indien.
802.11n-standarden fungerar på både 2,4 GHz- och 5,0 GHz-frekvenserna.
Detta gör att den kan vara bakåtkompatibel med 802.11a, 802.11b och 802.11g, förutsatt att basstationen har dubbla radioapparater.
Hastigheterna på 802.11n är betydligt snabbare än sina föregångare med en maximal teoretisk genomströmning på 600 Mbit/s.
Duvall, som är gift och har två vuxna barn, gjorde inget större intryck på Miller, som historien berättades för.
När han tillfrågades om en kommentar sa Miller: "Mike pratar mycket under utfrågningen... Jag gjorde mig i ordning så jag hörde inte riktigt vad han sa."
"Vi kommer att sträva efter att minska koldioxidutsläppen per BNP-enhet med en anmärkningsvärd marginal till 2020 från 2005 års nivå", sade Hu.
Han angav ingen siffra för nedskärningarna, utan sa att de kommer att göras baserat på Kinas ekonomiska produktion.
Hu uppmuntrade utvecklingsländerna "att undvika den gamla vägen att först förorena och sedan städa upp".
Han tillade att "de dock inte bör bli ombedda att ta på sig skyldigheter som går utöver deras utvecklingsstadium, ansvar och förmåga".
Iraq Study Group presenterade sin rapport klockan 12.00 GMT idag.
Den varnar för att ingen kan garantera att något agerande i Irak i nuläget kommer att stoppa sekteristisk krigföring, växande våld eller en glidning mot kaos.
Rapporten inleds med en vädjan om en öppen debatt och bildandet av ett samförstånd i USA om politiken gentemot Mellanöstern.
Betänkandet är mycket kritiskt till nästan varje aspekt av den verkställande maktens nuvarande politik gentemot Irak och uppmanar till en omedelbar kursändring.
Den första av de 78 rekommendationerna är att ett nytt diplomatiskt initiativ bör tas före årets slut för att säkra Iraks gränser mot fientliga ingripanden och för att återupprätta diplomatiska förbindelser med sina grannar.
Den nuvarande senatorn och argentinska första damen Cristina Fernández de Kirchner tillkännagav sin presidentkandidatur i går kväll i La Plata, en stad 50 kilometer från Buenos Aires.
Kirchner tillkännagav sin avsikt att kandidera till presidentposten på den argentinska teatern, samma plats som hon använde för att starta sin kampanj för senaten 2005 som medlem av Buenos Aires-provinsens delegation.
Debatten utlöstes av kontroverser om utgifter för katastrofhjälp och återuppbyggnad i kölvattnet av orkanen Katrina. som vissa finanspolitiskt konservativa skämtsamt har kallat "Bushs New Orleans-avtal".
Liberal kritik av återuppbyggnadsarbetet har fokuserat på tilldelningen av återuppbyggnadskontrakt till vad som uppfattas som Washingtons insiders.
Över fyra miljoner människor reste till Rom för att delta i begravningen.
Antalet närvarande var så stort att det inte var möjligt för alla att få tillträde till begravningen på Petersplatsen.
Flera stora tv-skärmar installerades på olika platser i Rom för att låta folket titta på ceremonin.
I många andra städer i Italien och i resten av världen, särskilt i Polen, gjordes liknande uppställningar, som sågs av ett stort antal människor.
Historiker har kritiserat tidigare FBI-policyer för att fokusera resurser på fall som är lätta att lösa, särskilt fall med stulna bilar, i syfte att öka byråns framgångsgrad.
Kongressen började finansiera obscenitetsinitiativet under budgetåret 2005 och specificerade att FBI måste ägna 10 agenter åt vuxenpornografi.
Robin Uthappa gjorde innings högsta poäng, 70 runs på bara 41 bollar genom att slå 11 fyror och 2 sexor.
Slagmännen Sachin Tendulkar och Rahul Dravid presterade bra och gjorde ett partnerskap på hundra runs.
Men efter att ha förlorat kaptenens wicket gjorde Indien bara 36 runs och förlorade 7 wickets för att avsluta innings.
USA:s president George W. Bush anlände till Singapore på morgonen den 16 november och inledde en veckolång rundresa i Asien.
Han hälsades välkommen av Singapores vice premiärminister Wong Kan Seng och diskuterade handels- och terrorismfrågor med Singapores premiärminister Lee Hsien Loong.
Efter en vecka av förluster i mellanårsvalet berättade Bush för en publik om den expanderande handeln i Asien.
Premiärminister Stephen Harper har gått med på att skicka regeringens "Clean Air Act" till en kommitté med alla partier för granskning, före dess andra behandling, efter tisdagens 25 minuter långa möte med NDP-ledaren Jack Layton vid PMO.
Layton hade bett om ändringar i de konservativas miljöproposition under mötet med premiärministern och bett om en "grundlig och fullständig omskrivning" av det konservativa partiets miljölag.
Ända sedan den federala regeringen gick in för att ta över finansieringen av Mersey-sjukhuset i Devonport, Tasmanien, har delstatsregeringen och vissa federala parlamentsledamöter kritiserat denna handling som ett jippo i förspelet till det federala valet som ska utlysas i november.
Men premiärminister John Howard har sagt att lagen bara var för att skydda sjukhusets faciliteter från att nedgraderas av den tasmanska regeringen, genom att ge ytterligare 45 miljoner australiska dollar.
Enligt den senaste bulletinen indikerade havsnivåmätningar att en tsunami genererades. Det fanns en viss tydlig tsunamiaktivitet i närheten av Pago Pago och Niue.
Inga större skador eller personskador har rapporterats i Tonga, men strömmen bröts tillfälligt, vilket enligt uppgift hindrade de tonganska myndigheterna från att ta emot tsunamivarningen som utfärdats av PTWC.
Fjorton skolor på Hawaii som ligger vid eller nära kusten var stängda hela onsdagen trots att varningarna hade hävts.
USA:s president George W. Bush välkomnade beskedet.
Bushs talesman Gordon Johndroe kallade Nordkoreas löfte "ett stort steg mot målet att uppnå en verifierbar kärnvapennedrustning på Koreahalvön".
Den tionde namngivna stormen under den atlantiska orkansäsongen, den subtropiska stormen Jerry, bildades i Atlanten idag.
National Hurricane Center (NHC) säger att Jerry i nuläget inte utgör något hot mot land.
U.S. Corps of Engineers uppskattade att 6 tum nederbörd skulle kunna bryta igenom de tidigare skadade vallarna.
Det nionde distriktet, som drabbades av översvämningar så högt som 20 meter under orkanen Katrina, ligger för närvarande i midjehögt vatten eftersom den närliggande fördämningen översvämmades.
Vatten rinner över vallen i en sektion som är 100 fot bred.
Commons administratör Adam Cuerden uttryckte sin frustration över raderingarna när han talade med Wikinews förra månaden.
"Han (Wales) ljög i princip för oss från början. För det första genom att agera som om detta var av juridiska skäl. För det andra genom att låtsas att han lyssnade på oss, ända fram till att han raderade sin konst."
Irritationen i samhället ledde till att man nu försöker utarbeta en policy för sexuellt innehåll för webbplatsen, som är värd för miljontals öppet licensierade medier.
Arbetet som utfördes var mestadels teoretiskt, men programmet skrevs för att simulera observationer gjorda av Skytten.
Effekten som teamet letade efter skulle orsakas av tidvattenkrafter mellan galaxens mörka materia och Vintergatans mörka materia.
Precis som månen utövar en dragningskraft på jorden och orsakar tidvatten, så utövar Vintergatan en kraft på Skyttens galax.
Forskarna kunde dra slutsatsen att den mörka materian påverkar annan mörk materia på samma sätt som vanlig materia gör.
Denna teori säger att den mesta mörka materian runt en galax finns runt en galax i en slags halo, och består av massor av små partiklar.
Tv-rapporter visar vit rök som kommer från anläggningen.
Lokala myndigheter varnar boende i närheten av anläggningen att stanna inomhus, stänga av luftkonditioneringen och inte dricka kranvatten.
Enligt Japans kärnkraftsmyndighet har radioaktivt cesium och jod identifierats vid anläggningen.
Myndigheterna spekulerar i att detta tyder på att behållare med uranbränsle på platsen kan ha spruckit och läcker.
Dr. Tony Moll upptäckte den extremt läkemedelsresistenta tuberkulosen (XDR-TB) i den sydafrikanska regionen KwaZulu-Natal.
I en intervju sa han att den nya varianten var "mycket oroande och alarmerande på grund av den mycket höga dödligheten".
En del patienter kan ha smittats på sjukhuset, tror dr Moll, och minst två av dem var sjukvårdspersonal på sjukhuset.
Under ett år kan en smittad person smitta 10–15 närkontakter.
Andelen XDR-TB i hela gruppen personer med tuberkulos verkar dock fortfarande vara låg. 6 000 av de totalt 330 000 personer som smittats vid en viss tidpunkt i Sydafrika.
Satelliterna, som båda vägde över 1 000 pund och färdades i cirka 17 500 miles per timme, kolliderade 491 miles ovanför jorden.
Forskare säger att explosionen som orsakades av kollisionen var massiv.
De försöker fortfarande avgöra hur stor kraschen var och hur jorden kommer att påverkas.
USA:s strategiska kommando vid det amerikanska försvarsdepartementets kontor spårar vrakdelarna.
Resultatet av plottningsanalysen kommer att publiceras på en offentlig webbplats.
En läkare som arbetade på Children's Hospital of Pittsburgh, Pennsylvania kommer att åtalas för grovt mord efter att hennes mamma hittades död i bagageutrymmet på sin bil i onsdags, säger myndigheterna i Ohio.
Dr. Malar Balasubramanian, 29, hittades i Blue Ash, Ohio, en förort cirka 15 mil norr om Cincinnati liggande på marken bredvid vägen i en T-shirt och underkläder i ett till synes tungt medicinerat tillstånd.
Hon dirigerade poliserna till sin svarta Oldsmobile Intrigue som låg 500 meter bort.
Där hittade de kroppen av Saroja Balasubramanian, 53, täckt av blodfläckade filtar.
Polisen sa att kroppen verkade ha legat där i ungefär ett dygn.
De första sjukdomsfallen den här säsongen rapporterades i slutet av juli.
Sjukdomen bärs av grisar, som sedan migrerar till människor via myggor.
Utbrottet har fått den indiska regeringen att vidta åtgärder som att placera ut grisfångare i hårt drabbade områden, dela ut tusentals mygggardiner och spruta bekämpningsmedel.
Regeringen har också utlovat flera miljoner flaskor med hjärninflammationsvaccin, vilket kommer att hjälpa till att förbereda hälsomyndigheterna för nästa år.
Planerna på att vaccin skulle levereras till de historiskt sett värst drabbade områdena i år försenades på grund av brist på pengar och låg prioritering i förhållande till andra sjukdomar.
1956 flyttade Słania till Sverige, där han tre år senare började arbeta för Posten och blev deras chefsgravör.
Han producerade över 1 000 frimärken för Sverige och 28 andra länder.
Hans arbete är av sådan erkänd kvalitet och detaljrikedom att han är ett av de mycket få "kända namnen" bland filatelisterna. Vissa specialiserar sig på att samla hans verk på egen hand.
Hans 1 000:e frimärke var den magnifika "Great Deeds by Swedish Kings" av David Klöcker Ehrenstrahl år 2000, som finns med i Guinness rekordbok.
Han var också engagerad i att gravera sedlar för många länder, bland annat porträtten av premiärministern på framsidan av de nya kanadensiska 5- och 100-dollarsedlarna.
Efter olyckan transporterades Gibson till sjukhus men avled kort därefter.
Lastbilschauffören, som är 64 år, skadades inte i kraschen.
Själva fordonet fördes bort från olycksplatsen cirka klockan 1200 GMT samma dag.
En person som arbetade i en bilverkstad i närheten av den plats där olyckan inträffade sade: "Det fanns barn som väntade på att få korsa vägen och alla skrek och grät."
De sprang alla tillbaka från platsen där olyckan hade inträffat.
Andra frågor som står på dagordningen på Bali är att rädda världens återstående skogar och dela med sig av teknik för att hjälpa utvecklingsländer att växa på mindre förorenande sätt.
FN hoppas också kunna färdigställa en fond för att hjälpa länder som drabbats av den globala uppvärmningen att hantera effekterna.
Pengarna skulle kunna gå till översvämningssäkra hus, bättre vattenhantering och diversifiering av grödor.
Fluke skrev att vissa försök att överrösta kvinnor från att tala ut om kvinnors hälsa misslyckades.
Hon kom fram till denna slutsats på grund av de många positiva kommentarer och uppmuntran som skickades till henne från både kvinnliga och manliga individer som uppmanade till att preventivmedel skulle betraktas som en medicinsk nödvändighet.
När striderna upphörde efter att de sårade transporterats till sjukhuset stannade ett 40-tal av de andra fångarna kvar på gården och vägrade återvända till sina celler.
Förhandlarna försökte rätta till situationen, men fångarnas krav är oklara.
Mellan 22:00-23:00 MDT startades en brand av de intagna på gården.
Snart kom kravallutrustade poliser in på gården och trängde in fångarna i ett hörn med tårgas.
Räddningstjänsten släckte till slut branden vid 23.35-tiden.
Efter att dammen byggdes 1963 stoppades de säsongsbetonade översvämningarna som skulle sprida sediment i hela floden.
Detta sediment var nödvändigt för att skapa sandbankar och stränder, som fungerade som livsmiljöer för vilda djur.
Som ett resultat av detta har två fiskarter dött ut och två andra har blivit utrotningshotade, däribland knölfärnan.
Även om vattennivån bara kommer att stiga några meter efter översvämningen, hoppas myndigheterna att det kommer att räcka för att återställa eroderade sandbankar nedströms.
Ingen tsunamivarning har utfärdats, och enligt Jakartas geofysiska byrå kommer ingen tsunamivarning att utfärdas eftersom skalvet inte uppfyllde kravet på magnituden 6,5.
Trots att det inte fanns något tsunamihot började invånarna få panik och började lämna sina företag och hem.
Även om Winfrey var tårögd i sitt avsked gjorde hon det klart för sina fans att hon kommer tillbaka.
"Det här kommer inte att bli ett farväl. Detta är slutet på ett kapitel och början på ett nytt."
Slutresultatet från president- och parlamentsvalen i Namibia har visat att den sittande presidenten Hifikepunye Pohamba har blivit omvald med stor marginal.
Det styrande partiet, South West Africa People's Organisation (SWAPO), behöll också majoriteten i parlamentsvalet.
Koalitionstrupper och afghanska trupper har gått in i området för att säkra platsen och andra koalitionsflygplan har skickats för att hjälpa till.
Kraschen inträffade högt upp i bergig terräng och tros ha varit resultatet av fientlig eld.
Arbetet med att söka efter nedslagsplatsen möts av dåligt väder och tuff terräng.
Den medicinska välgörenhetsorganisationen Mangola, Läkare utan gränser och Världshälsoorganisationen WHO säger att det är det värsta utbrottet som registrerats i landet.
Richard Veerman, talesman för Läkare utan gränser, sade: "Angola är på väg mot sitt värsta utbrott någonsin och situationen är fortfarande mycket dålig i Angola", sade han.
Matcherna startade klockan 10:00 med bra väder och bortsett från duggregn på förmiddagen som snabbt klarnade upp var det en perfekt dag för 7:s rugby.
Turneringens toppseedade Sydafrika började på rätt sätt när de vann komfortabelt med 26–00 mot 5:e-seedade Zambia.
Sydafrika såg klart ringrostiga ut i matchen mot sina sydliga systrar, men förbättrades stadigt allt eftersom turneringen fortskred.
Deras disciplinerade försvar, bollbehandling och utmärkta lagarbete gjorde att de stack ut och det var tydligt att detta var laget att slå.
Tjänstemän för staden Amsterdam och Anne Frank-museet uppger att trädet är infekterat med en svamp och utgör en folkhälsorisk eftersom de hävdar att det var i överhängande fara att falla omkull.
Den skulle ha klippts ner på tisdagen, men räddades efter ett nöddomstolsbeslut.
Alla grottöppningar, som fick namnet "De sju systrarna", är minst 100 till 250 meter (328 till 820 fot) i diameter.
Infraröda bilder visar att temperaturvariationerna från natt och dag visar att det sannolikt rör sig om grottor.
– De är svalare än den omgivande ytan på dagen och varmare på natten.
Deras termiska beteende är inte lika stabilt som stora grottor på jorden som ofta håller en ganska konstant temperatur, men det stämmer överens med att dessa är djupa hål i marken, säger Glen Cushing från United States Geological Survey (USGS) Astrogeology Team och Northern Arizona University i Flagstaff, Arizona.
I Frankrike har röstning traditionellt sett varit en lågteknologisk upplevelse: väljarna isolerar sig i ett bås och lägger ett förtryckt pappersark som anger vilken kandidat de vill rösta på i ett kuvert.
Efter att tjänstemännen har verifierat väljarens identitet lägger väljaren kuvertet i valurnan och undertecknar röstlängden.
Den franska vallagen är ganska strikt kodifierad av förfarandet.
Sedan 1988 måste valurnorna vara genomskinliga så att väljare och observatörer kan intyga att det inte finns några kuvert när omröstningen inleds och att inga kuvert läggs till förutom de som tillhör de vederbörligen räknade och behöriga väljarna.
Kandidater kan skicka representanter för att bevittna varje del av processen. På kvällen räknas rösterna av volontärer under hård övervakning, enligt särskilda procedurer.
ASUS Eee PC, som tidigare lanserats över hela världen för kostnadsbesparing och funktionalitetsfaktorer, blev ett hett ämne under Taipei IT Month 2007.
Men konsumentmarknaden för bärbara datorer kommer att bli radikalt varierad och förändrad efter att ASUS tilldelades 2007 års Taiwan Sustainable Award av Executive Yuan i Republiken Kina.
På stationens hemsida beskrivs showen som "old school radio theatre with a new and outrageous geeky twist!"
I början visades programmet enbart på den långvariga internetradiosajten TogiNet Radio, en webbplats som fokuserade på pratradio.
I slutet av 2015 etablerade TogiNet AstroNet Radio som en dotterstation.
Serien hade ursprungligen amatörröstskådespelare från östra Texas.
Den utbredda plundringen ska ha fortsatt under natten, eftersom poliser inte var närvarande på Bisjkeks gator.
Bisjkek beskrevs som på väg in i ett tillstånd av "anarki" av en observatör, då gäng av människor strövade omkring på gatorna och plundrade butiker på konsumtionsvaror.
Flera invånare i Bisjkek beskyllde demonstranter från söder för laglösheten.
Sydafrika har besegrat All Blacks (Nya Zeeland) i en rugby union Tri Nations match på Royal Bafokeng Stadium i Rustenburg, Sydafrika.
Slutresultatet blev en enpoängsseger, 21 mot 20, vilket avslutade All Blacks 15 matcher långa segersvit.
För Springboks innebar det slutet på en fem matcher lång förlustsvit.
Det var den sista matchen för All Blacks, som redan hade vunnit trofén för två veckor sedan.
Den sista matchen i serien kommer att äga rum på Ellis Park i Johannesburg nästa vecka, när Springboks spelar mot Australien.
En måttlig jordbävning skakade västra Montana klockan 22.08 på måndagen.
Inga omedelbara rapporter om skador har mottagits av United States Geological Survey (USGS) och dess National Earthquake Information Center.
Jordbävningen hade sitt centrum omkring 20 km nord-nordost om Dillon och omkring 65 km söder om Butte.
Den för människor dödliga fågelinfluensastammen, H5N1, har bekräftats ha smittat en död vildand som hittades i måndags i ett träsk nära Lyon i östra Frankrike.
Frankrike är det sjunde landet i EU som drabbats av detta virus. Österrike, Tyskland, Slovenien, Bulgarien, Grekland och Italien.
Misstänkta fall av H5N1 i Kroatien och Danmark är fortfarande obekräftade.
Chambers hade stämt Gud för "utbredd död, förstörelse och terrorisering av miljoner och åter miljoner av jordens invånare".
Chambers, som är agnostiker, hävdar att hans stämningsansökan är "oseriös" och att "vem som helst kan stämma vem som helst".
Berättelsen som presenteras i den franska operan, av Camille Saint-Saëns, handlar om en konstnär "vars liv dikteras av en kärlek till droger och Japan".
Som ett resultat av detta röker artisterna cannabisjointar på scenen, och teatern själv uppmuntrar publiken att delta.
Den tidigare talmannen i representanthuset Newt Gingrich, Texas guvernör Rick Perry och kongressledamoten Michele Bachmann slutade på fjärde, femte respektive sjätte plats.
Efter att resultaten kommit in hyllade Gingrich Santorum, men hade hårda ord för Romney, på vars vägnar negativa kampanjannonser sändes i Iowa mot Gingrich.
Perry uppgav att han skulle "återvända till Texas för att utvärdera resultaten av kvällens caucus, avgöra om det finns en väg framåt för mig själv i det här loppet", men sa senare att han skulle stanna kvar i tävlingen och tävla i primärvalet i South Carolina den 21 januari.
Bachmann, som vann Ames Straw Poll i augusti, bestämde sig för att avsluta sin kampanj.
Fotografen transporterades till Ronald Reagan UCLA Medical Center, där han senare avled.
Han ska ha varit i 20-årsåldern. I ett uttalande sa Bieber: "Även om jag inte var närvarande eller direkt involverad i denna tragiska olycka, är mina tankar och böner med offrets familj."
Nöjesnyhetssajten TMZ förstår att fotografen stannade sitt fordon på andra sidan Sepulveda Boulevard och försökte ta bilder av polisstoppet innan han korsade vägen och fortsatte, vilket fick California Highway Patrol-polisen som genomförde trafikstoppet att beordra honom tillbaka över, två gånger.
Enligt polisen är det osannolikt att föraren av fordonet som körde på fotografen kommer att åtalas.
Med endast arton medaljer tillgängliga per dag har ett antal länder misslyckats med att ta sig upp på medaljpallen.
Bland dem finns Nederländerna, där Anna Jochemsen slutade på nionde plats i damernas stående klass i super-G i går, och Finland där Katja Saarinen slutade på tionde plats i samma tävling.
Australiens Mitchell Gourley slutade på elfte plats i herrarnas stående Super-G. Tjecken Oldrich Jelinek slutade på sextonde plats i herrarnas sittande super-G.
Arly Velasquez från Mexiko slutade på femtonde plats i herrarnas sittande super-G. Nya Zeelands Adam Hall slutade på nionde plats i herrarnas stående Super-G.
Polens synskadade skidåkare Maciej Krezel och guiden Anna Ogarzynska slutade på trettonde plats i super-G. Sydkoreas Jong Seork Park slutade på tjugofjärde plats i herrarnas sittande super-G.
FN:s fredsbevarande styrkor, som anlände till Haiti efter jordbävningen 2010, beskylls för spridningen av sjukdomen som började nära truppernas läger.
Enligt stämningsansökan desinficerades inte avfallet från FN-lägret ordentligt, vilket ledde till att bakterier kom in i bifloden Artibonite, en av Haitis största.
Innan trupperna anlände hade Haiti inte stött på problem relaterade till sjukdomen sedan 1800-talet.
Haitiska institutet för rättvisa och demokrati har hänvisat till oberoende studier som tyder på att den nepalesiska FN:s fredsbevarande bataljon ovetandes förde sjukdomen till Haiti.
Danielle Lantagne, FN:s expert på sjukdomen, uppgav att utbrottet troligen orsakades av de fredsbevarande styrkorna.
Hamilton bekräftade att Howard University Hospital tog emot patienten i stabilt tillstånd.
Patienten hade varit i Nigeria, där några fall av ebolaviruset har förekommit.
Sjukhuset har följt protokoll för infektionskontroll, inklusive att separera patienten från andra för att förhindra eventuell infektion av andra.
Innan The Simpsons hade Simon arbetat med flera serier i olika positioner.
Under 1980-talet arbetade han med program som Taxi, Cheers och The Tracy Ullman Show.
1989 hjälpte han till att skapa The Simpsons tillsammans med Brooks och Groening, och var ansvarig för att anställa seriens första manusteam.
Trots att han lämnade serien 1993 behöll han titeln som exekutiv producent och fortsatte att få tiotals miljoner dollar varje säsong i royalties.
Tidigare rapporterade den kinesiska nyhetsbyrån Xinhua att ett plan kapats.
Senare rapporter uppgav att planet mottog ett bombhot och omdirigerades tillbaka till Afghanistan och landade i Kandahar.
De tidiga rapporterna säger att planet omdirigerades tillbaka till Afghanistan efter att ha nekats en nödlandning i Ürümqi.
Flygolyckor är vanliga i Iran, som har en åldrande flotta som är dåligt underhållen både för civila och militära operationer.
Internationella sanktioner har inneburit att nya flygplan inte kan köpas.
Tidigare i veckan kraschade en polishelikopter som dödade tre personer och skadade ytterligare tre.
Förra månaden drabbades Iran av sin värsta flygkatastrof på flera år när ett flygplan på väg till Armenien kraschade och de 168 ombord omkom.
Samma månad körde ett annat flygplan över en landningsbana i Mashhad och kolliderade med en vägg och dödade sjutton personer.
Aerosmith har ställt in sina återstående konserter på sin turné.
Rockbandet skulle turnera i USA och Kanada fram till den 16 september.
De har ställt in turnén efter att sångaren Steven Tyler skadades efter att han föll av scenen när han uppträdde den 5 augusti.
Murray förlorade första set i tiebreak efter att båda männen hållit varsin serve i setet.
Del Potro hade ett tidigt övertag i andra set, men även detta krävde ett tiebreak efter att ha nått 6-6.
Potro fick behandling för sin axel vid denna tidpunkt men lyckades återvända till matchen.
Programmet startade klockan 20.30 lokal tid (15.00 UTC).
Kända sångare över hela landet framförde bhajans, eller hängivna sånger, till Shri Shyams fötter.
Sångaren Sanju Sharma inledde kvällen, följd av Jai Shankar Choudhary. Esented Chhappan bhog bhajan också. Sångaren Raju Khandelwal ackompanjerade honom.
Sedan tog Lakkha Singh ledningen i att sjunga bhajans.
108 tallrikar med Chhappan Bhog (inom hinduismen 56 olika ätbara föremål, som godis, frukt, nötter, rätter etc. som offras till gudomen) serverades till Baba Shyam.
Lakkha Singh presenterade också chhappan bhog bhajan. Sångaren Raju Khandelwal ackompanjerade honom.
Vid torsdagens keynote-presentation av Tokyo Game Show avslöjade Nintendos president Satoru Iwata kontrollerdesignen för företagets nya Nintendo Revolution-konsol.
Styrenheten liknar en TV-fjärrkontroll och använder två sensorer placerade nära användarens TV för att triangulera dess position i tredimensionellt utrymme.
Detta gör det möjligt för spelare att styra handlingar och rörelser i videospel genom att flytta enheten genom luften.
Giancarlo Fisichella tappade kontrollen över sin bil och avslutade loppet mycket snart efter starten.
Hans teamkamrat Fernando Alonso var i ledningen under större delen av loppet, men bröt det direkt efter sitt depåstopp, förmodligen på grund av ett dåligt instucket höger framhjul.
Michael Schumacher avslutade sitt lopp inte långt efter Alonso, på grund av fjädringsskadorna i de många striderna under loppet.
"Hon är väldigt söt och sjunger ganska bra också", sa han enligt en utskrift av presskonferensen.
"Jag blev rörd varje gång vi repeterade om det här, från djupet av mitt hjärta."
Cirka 3 minuter in i uppskjutningen visade en inbyggd kamera att många bitar av isoleringsskum lossnade från bränsletanken.
De tros dock inte ha orsakat några skador på skytteln.
NASA:s chef för rymdfärjeprogrammet, N. Wayne Hale Jr., sade att skummet hade fallit "efter den tid vi är oroliga för".
Fem minuter in i displayen börjar en vind rulla in, ungefär en minut senare når vinden 70 km/h... Sen kommer regnet, men så hårt och så stort att det slår mot huden som en nål, sedan föll hagel från himlen, folk som fick panik och skrek och körde över varandra.
Jag förlorade min syster och hennes vän, och på vägen dit var det två funktionshindrade personer i rullstol, människor som bara hoppade över och knuffade dem, säger Armand Versace.
NHK rapporterade också att kärnkraftverket Kashiwazaki Kariwa i Niigata-prefekturen fungerade normalt.
Hokuriku Electric Power Co. rapporterade inga effekter av jordbävningen och att reaktor nummer 1 och 2 vid kärnkraftverket Shika stängdes.
Det rapporteras att cirka 9400 hushåll i regionen är utan vatten och cirka 100 utan el.
Vissa vägar har skadats, järnvägstrafiken har avbrutits i de drabbade områdena och flygplatsen Noto i prefekturen Ishikawa är fortfarande stängd.
En bomb exploderade utanför generalguvernörens kontor.
Ytterligare tre bomber exploderade nära regeringsbyggnader under loppet av två timmar.
Vissa rapporter anger den officiella dödssiffran till åtta, och officiella rapporter bekräftar att upp till 30 skadades. Men de slutliga siffrorna är ännu inte kända.
Både cyanursyra och melamin hittades i urinprover från husdjur som dött efter att ha ätit förorenat djurfoder.
De två föreningarna reagerar med varandra för att bilda kristaller som kan blockera njurfunktionen, säger forskare vid universitetet.
Forskarna observerade kristaller som bildades i katturin genom tillsats av melamin och cyanursyra.
Sammansättningen av dessa kristaller matchar de som finns i urinen hos drabbade husdjur jämfört med infraröd spektroskopi (FTIR).
Jag vet inte om du inser det eller inte, men de flesta varor från Centralamerika kom in i landet tullfritt.
Ändå beskattades åttio procent av våra varor genom tullar i de centralamerikanska länderna. Vi behandlar dig.
Det verkade inte vettigt för mig; Det var verkligen inte rättvist.
Allt jag säger till människor är att ni behandlar oss som vi behandlar er.
Kaliforniens guvernör Arnold Schwarzenegger undertecknade ett lagförslag som förbjuder försäljning eller uthyrning av våldsamma videospel till minderåriga.
Lagförslaget kräver att våldsamma videospel som säljs i delstaten Kalifornien ska märkas med en dekal med texten "18" och gör att försäljning till en minderårig straffas med böter på 1000 dollar per brott.
Riksåklagaren, Kier Starmer QC, gjorde ett uttalande i morse där han meddelade att både Huhne och Pryce åtalas.
Huhne har avgått och han kommer att ersättas i kabinettet av parlamentsledamoten Ed Davey. Parlamentsledamoten Norman Lamb förväntas ta över jobbet som näringsminister som Davey lämnar.
Huhne och Pryce ska infinna sig i Westminster Magistrates Court den 16 februari.
De omkomna var Nicholas Alden, 25, och Zachary Cuddeback, 21. Cuddeback hade varit chaufför.
Edgar Veguilla fick sår i armar och käkar medan Kristoffer Schneider fick genomgå rekonstruktiv kirurgi i ansiktet.
Ukas vapen misslyckades när det riktades mot en femte mans huvud. Schneider har pågående smärta, blindhet på ena ögat, en saknad del av skallen och ett ansikte som byggts om av titan.
Schneider vittnade via videolänk från en USAF-bas i sitt hemland.
Utöver onsdagens tävling tävlade Carpanedo i två individuella lopp i mästerskapen.
Hennes första var slalom, där hon fick en Not Finish i sitt första åk. 36 av de 116 tävlande hade samma resultat i det loppet.
I hennes andra tävling, storslalom, slutade hon på tionde plats i damernas sittgrupp med en sammanlagd tid på 4:41.30, 2:11.60 minuter långsammare än österrikiskan Claudia Loesch och 1:09.02 minuter långsammare än Gyöngyi Dani från Ungern som slutade på nionde plats.
Fyra åkare i damernas sittgrupp misslyckades med att fullfölja sina åk, och 45 av de totalt 117 åkarna i storslalom misslyckades med att placera sig i loppet.
Polisen i Madhya Pradesh återfann den stulna bärbara datorn och mobiltelefonen.
Biträdande generalinspektör D K Arya sa: "Vi har gripit fem personer som våldtog den schweiziska kvinnan och återtog hennes mobil och bärbara dator".
De anklagade heter Baba Kanjar, Bhutha Kanjar, Rampro Kanjar, Gaza Kanjar och Vishnu Kanjar.
Polisinspektör Chandra Shekhar Solanki sade att de anklagade dök upp i rätten med täckta ansikten.
Trots att tre personer befann sig i huset när bilen kolliderade med det, skadades ingen av dem.
Föraren fick dock allvarliga skador i huvudet.
Vägen där olyckan inträffade stängdes tillfälligt av medan räddningstjänsten befriade föraren från den röda Audi TT.
Han var först inlagd på James Paget Hospital i Great Yarmouth.
Han flyttades därefter till Addenbrooke's Hospital i Cambridge.
Adekoya har sedan dess suttit i Edinburgh Sheriff Court anklagad för att ha mördat sin son.
Hon sitter häktad i väntan på åtal och rättegång, men eventuella ögonvittnesbevis kan vara befläckade eftersom hennes bild har fått stor spridning.
Detta är vanligt på andra håll i Storbritannien, men det skotska rättsväsendet fungerar annorlunda och domstolar har betraktat publicering av foton som potentiellt skadligt.
Professor Pamela Ferguson vid University of Dundee noterar att "journalister verkar gå på en farlig linje när de publicerar bilder etc av misstänkta".
Crown Office, som har det övergripande ansvaret för åtal, har meddelat journalister att inga ytterligare kommentarer kommer att ges åtminstone fram till åtalet.
Dokumentet kommer, enligt läckan, att hänvisa till gränstvisten, som Palestina vill ha baserat på gränserna före Mellanösternkriget 1967.
Andra ämnen som tas upp är enligt uppgift den framtida staten Jerusalem, som är helig för båda nationerna, och frågan om Jordandalen.
Israel kräver en fortsatt militär närvaro i dalen i tio år när ett avtal väl är undertecknat, medan den palestinska myndigheten går med på att bara lämna sådan närvaro i fem år.
Skyttarna i det kompletterande bekämpningsförsöket skulle övervakas noggrant av parkvakter, eftersom försöket övervakades och dess effektivitet utvärderades.
I ett samarbete mellan NPWS och Sporting Shooters Association of Australia (NSW) Inc rekryterades kvalificerade volontärer inom ramen för Sporting Shooters Associations jaktprogram.
Enligt Mick O'Flynn, tillförordnad chef för parkbevarande och kulturarv vid NPWS, fick de fyra skyttar som valdes ut för den första skjutoperationen omfattande säkerhets- och utbildningsinstruktioner.
Martelly svor i går in ett nytt provisoriskt valråd (CEP) med nio medlemmar.
Det är Martellys femte CEP på fyra år.
Förra månaden rekommenderade en presidentkommission den tidigare CEP:s avgång som en del av ett åtgärdspaket för att föra landet mot nyval.
Uppdraget var Martellys svar på de omfattande protesterna mot regimen som började i oktober.
De stundtals våldsamma protesterna utlöstes av att val inte hölls, varav vissa skulle ha hållits sedan 2011.
Omkring 60 fall av överhettning av iPod-enheter som inte fungerar som de ska har rapporterats, vilket har orsakat totalt sex bränder och lämnat fyra personer med mindre brännskador.
Japans ministerium för ekonomi, handel och industri (METI) sade att det hade varit medvetet om 27 olyckor relaterade till enheterna.
Förra veckan meddelade METI att Apple hade informerat dem om ytterligare 34 överhettningsincidenter, som företaget kallade "icke-allvarliga".
Departementet svarade med att kalla Apples uppskjutande av rapporten "verkligen beklagligt".
Jordbävningen drabbade Mariana klockan 07:19 lokal tid (21:19 GMT på fredagen).
Nordmarianernas krisledningskontor sade att det inte fanns några skador rapporterade i landet.
Även Pacific Tsunami Warning Center sade att det inte fanns någon indikation på tsunami.
En före detta filippinsk polis har hållit Hongkongs turister som gisslan genom att kapa deras buss i Filippinernas huvudstad Manila.
Rolando Mendoza avfyrade sitt M16-gevär mot turisterna.
Flera gisslan har räddats och minst sex har hittills bekräftats döda.
Sex personer som tagits som gisslan, däribland barn och äldre, släpptes i förtid, liksom de filippinska fotograferna.
Fotograferna tog senare en äldre dams plats när hon behövde toaletten. Mendoza sköts ner.
Liggins följde i sin fars fotspår och inledde en karriär inom medicin.
Han utbildade sig till förlossningsläkare och började arbeta på Aucklands National Women's Hospital 1959.
Medan han arbetade på sjukhuset började Liggins undersöka för tidig förlossning på sin fritid.
Hans forskning visade att om ett hormon administrerades skulle det påskynda fostrets lungmognad.
Xinhua rapporterade att regeringens utredare återfann två "svarta lådan" på onsdagen.
Andra brottare hyllade också Luna.
Tommy Dreamer sa: "Luna var den första drottningen av Extreme. Min första chef. Luna gick bort på natten av två månar. Ganska unik precis som hon. Stark kvinna."
Dustin "Goldust" Runnels kommenterade att "Luna var lika galen som jag... kanske till och med mer... älskar henne och kommer att sakna henne ... Förhoppningsvis är hon på en bättre plats."
Av 1 400 personer som tillfrågades inför det federala valet 2010 har de som motsätter sig att Australien blir en republik ökat med 8 procent sedan 2008.
Premiärministern Julia Gillard hävdade under kampanjen i det federala valet 2010 att hon ansåg att Australien skulle bli en republik i slutet av drottning Elizabeth II:s regeringstid.
34 procent av de tillfrågade delar denna uppfattning och vill att drottning Elizabeth II ska bli Australiens sista monark.
29 procent av de tillfrågade anser att Australien bör bli en republik så snart som möjligt, medan 31 procent anser att Australien aldrig bör bli en republik.
Den olympiska guldmedaljören skulle ha simmat i 100 och 200 meter frisim och i tre stafetter vid Samväldesspelen, men på grund av hans klagomål har hans kondition ifrågasatts.
Han har inte kunnat ta de droger som behövs för att övervinna sin smärta eftersom de är förbjudna från spelen.
Curtis Cooper, matematiker och professor i datavetenskap vid University of Central Missouri, upptäckte det största kända primtalet hittills den 25 januari.
Flera personer verifierade upptäckten med hjälp av olika hård- och mjukvara i början av februari och det tillkännagavs på tisdagen.
Kometer kan möjligen ha varit en källa till vattentillförsel till jorden tillsammans med organiskt material som kan bilda proteiner och stödja liv.
Forskare hoppas kunna förstå hur planeter bildas, särskilt hur jorden bildades, eftersom kometer kolliderade med jorden för länge sedan.
Cuomo, 53, började sin guvernörsperiod tidigare i år och undertecknade förra månaden ett lagförslag som legaliserar samkönade äktenskap.
Han refererade till ryktena som "politiskt prat och dumheter".
Det spekuleras i att han kommer att ställa upp i presidentvalet 2016.
NextGen är ett system som FAA hävdar skulle göra det möjligt för flygplan att flyga kortare rutter och spara miljontals liter bränsle varje år och minska koldioxidutsläppen.
Den använder satellitbaserad teknik i motsats till äldre markradarbaserad teknik för att göra det möjligt för flygledare att lokalisera flygplan med större precision och ge piloter mer exakt information.
Inga extra transporter sätts in och tåg ovan jord kommer inte att stanna vid Wembley, och parkering och infartsparkeringar är inte tillgängliga på marken.
Rädslan för brist på transporter gjorde att matchen skulle tvingas spelas bakom stängda dörrar utan lagets supportrar.
En studie som publicerades på torsdagen i tidskriften Science rapporterade om bildandet av en ny fågelart på de ecuadorianska Galápagosöarna.
Forskare från Princeton University i USA och Uppsala universitet i Sverige rapporterade att den nya arten utvecklades på bara två generationer, även om denna process har ansetts ta mycket längre tid, på grund av häckning mellan en endemisk darwinfink, Geospiza fortes, och den invandrade kaktusfinken, Geospiza conirostris.
Guld kan bearbetas till alla möjliga former. Den kan rullas till små former.
Den kan dras till tunn tråd, som kan vridas och flätas. Den kan hamras eller rullas till ark.
Den kan göras mycket tunn och fästas på annan metall. Den kan göras så tunn att den ibland användes för att dekorera de handmålade bilderna i böcker som kallas "illuminerade manuskript".
Detta kallas en kemikalies pH. Du kan göra en indikator med rödkålsjuice.
Kåljuicen ändrar färg beroende på hur sur eller basisk (alkalisk) kemikalien är.
pH-nivån indikeras av mängden vätejoner (H i pH) i den testade kemikalien.
Vätejoner är protoner som fick sina elektroner avskalade från dem (eftersom väteatomer består av en proton och en elektron).
Snurra ihop de två torra pulvren och pressa dem sedan till en boll med rena, våta händer.
Fukten på dina händer kommer att reagera med de yttre lagren, vilket kommer att kännas roligt och bilda ett slags skal.
Städerna Harappa och Mohenjo-daro hade en vattentoalett i nästan varje hus, ansluten till ett sofistikerat avloppssystem.
Rester av avloppssystem har hittats i husen i de minoiska städerna Kreta och Santorini i Grekland.
Det fanns också toaletter i forntida Egypten, Persien och Kina. I den romerska civilisationen var toaletter ibland en del av offentliga badhus där män och kvinnor var tillsammans i blandat sällskap.
När du ringer någon som är tusentals mil bort använder du en satellit.
Satelliten i rymden tar emot samtalet och reflekterar det sedan nedåt igen, nästan omedelbart.
Satelliten skickades ut i rymden med en raket. Forskare använder teleskop i rymden eftersom jordens atmosfär förvränger en del av vårt ljus och vår syn.
Det krävs en gigantisk raket som är över 100 meter hög för att placera en satellit eller ett teleskop i rymden.
Hjulet har förändrat världen på otroliga sätt. Det största som hjulet har gjort för oss är att det har gett oss mycket enklare och snabbare transporter.
Det har gett oss tåget, bilen och många andra transportmedel.
Under dem finns fler medelstora katter som äter medelstora byten, allt från kaniner till antiloper och rådjur.
Slutligen finns det många små katter (inklusive lösa sällskapskatter) som äter de mycket mer talrika små bytena som insekter, gnagare, ödlor och fåglar.
Hemligheten bakom deras framgång är konceptet med nischen, ett speciellt jobb som varje katt har och som hindrar den från att konkurrera med andra.
Lejon är de mest sociala katterna och lever i stora grupper som kallas flockar.
Flockar består av en till tre besläktade vuxna hanar, tillsammans med så många som trettio honor och ungar.
Honorna är vanligtvis nära släkt med varandra och är en stor familj av systrar och döttrar.
Lejonflockar beter sig ungefär som flockar av vargar eller hundar, djur som är förvånansvärt lika lejon (men inte andra stora kattdjur) i beteende, och som också är mycket dödliga för sina byten.
Tigern är en mångsidig atlet som kan klättra (men inte bra), simma, hoppa långa sträckor och dra med fem gånger kraften hos en stark människa.
Tigern tillhör samma grupp (Släkte Panthera) som lejon, leoparder och jaguarer. Dessa fyra katter är de enda som kan ryta.
Tigerns rytande är inte som ett lejons högljudda rytande, utan mer som en mening av snarkiga, skrikande ord.
Ozeloter gillar att äta smådjur. De kommer att fånga apor, ormar, gnagare och fåglar om de kan. Nästan alla djur som ozeloten jagar är mycket mindre än vad den är.
Forskare tror att ozeloter följer efter och hittar djur att äta (byten) genom lukten och sniffar efter var de har varit på marken.
De kan se mycket bra i mörker med mörkerseende och rör sig också mycket smygande. Ozeloter jagar sitt byte genom att smälta in i sin omgivning och sedan kasta sig över sitt byte.
När en liten grupp levande varelser (en liten population) separeras från huvudpopulationen som de kom från (som om de flyttar över en bergskedja eller en flod, eller om de flyttar till en ny ö så att de inte lätt kan flytta tillbaka) kommer de ofta att befinna sig i en annan miljö än de var i tidigare.
Denna nya miljö har andra resurser och olika konkurrenter, så den nya befolkningen kommer att behöva andra funktioner eller anpassningar för att vara en stark konkurrent än vad de hade behövt tidigare.
Den ursprungliga populationen har inte förändrats alls, de behöver fortfarande samma anpassningar som tidigare.
Med tiden, när den nya populationen börjar anpassa sig till sin nya miljö, börjar de se mindre och mindre ut som den andra populationen.
Så småningom, efter tusentals eller till och med miljontals år, kommer de två populationerna att se så olika ut att de inte kan kallas samma art.
Vi kallar denna process för artbildning, vilket helt enkelt betyder bildandet av nya arter. Artbildning är en oundviklig konsekvens och en mycket viktig del av evolutionen.
Växter producerar syre som människor andas, och de tar upp koldioxid som människor andas ut (det vill säga andas ut).
Växter får sin föda från solen genom fotosyntes. De ger också skugga.
Vi gör våra hus av växter och kläder av växter. De flesta livsmedel som vi äter är växter. Utan växter skulle djuren inte kunna överleva.
Mosasaurus var sin tids toppredatorer, så den fruktade ingenting, förutom andra mosasaurier.
Dess långa käkar var översållade med mer än 70 rakbladsvassa tänder, tillsammans med en extra uppsättning i gommen, vilket innebar att det inte fanns någon flyktväg för något som korsade dess väg.
Vi vet inte säkert, men den kan ha haft en kluven tunga. Dess föda bestod av sköldpaddor, stora fiskar, andra mosasaurier, och den kan till och med ha varit en kannibal.
Den attackerade också allt som kom in i vattnet; Inte ens en gigantisk dinosaurie som T. rex skulle vara någon match för den.
Även om det mesta av deras mat skulle vara bekant för oss, hade romarna sin beskärda del av konstiga eller ovanliga festföremål, inklusive vildsvin, påfågel, sniglar och en typ av gnagare som kallas hasselmus
En annan skillnad var att medan de fattiga och kvinnan åt sin mat sittande i stolar, tyckte de rika männen om att ha banketter tillsammans där de slappnade av på sidan medan de åt sina måltider.
Forntida romerska måltider kan inte ha inkluderat mat som kom till Europa från Amerika eller från Asien under senare århundraden.
De hade till exempel varken majs, tomater, potatis eller kakao, och ingen forntida romare smakade någonsin på en kalkon.
Babylonierna byggde var och en av sina gudar ett primärt tempel som ansågs vara gudens hem.
Folk offrade till gudarna och prästerna försökte tillgodose gudarnas behov genom ceremonier och festivaler.
Varje tempel hade en öppen tempelgård och sedan en inre helgedom som bara prästerna kunde gå in i.
Ibland byggdes speciella pyramidformade torn, så kallade ziggurater, för att vara en del av templen.
Toppen av tornet var en särskild helgedom för guden.
I det varma klimatet i Mellanöstern var huset inte så viktigt.
Det mesta av den hebreiska familjens liv ägde rum under bar himmel.
Kvinnorna lagade mat på gården; Butikerna var bara öppna diskar som vette ut mot gatan. Sten användes för att bygga hus.
Det fanns inga stora skogar i Kanaans land, så virke var mycket dyrt.
Grönland var glest befolkat. I de nordiska sagorna sägs det att Erik den Röde blev landsförvisad från Island för mord, och när han reste längre västerut hittade han Grönland och gav det namnet Grönland.
Men oavsett hans upptäckt bodde eskimåstammar redan där vid den tiden.
Även om varje land var "skandinaviskt" fanns det många skillnader mellan folket, kungarna, sederna och historien i Danmark, Sverige, Norge och Island.
Om du har sett filmen National Treasure kanske du tror att en skattkarta skrevs på baksidan av självständighetsförklaringen.
Det är dock inte sant. Även om det står något på baksidan av dokumentet är det inte en skattkarta.
På baksidan av självständighetsförklaringen stod det "Original Declaration of Independence daterad 4 juli 1776". Texten visas upp och ned längst ned i dokumentet.
Även om ingen med säkerhet vet vem som skrev det, är det känt att tidigt i dess liv rullades det stora pergamentdokumentet (det mäter 293/4 tum gånger 241/2 tum) ihop för förvaring.
Så det är troligt att notationen lades till helt enkelt som en etikett.
Landstigningarna på D-dagen och de följande striderna hade befriat norra Frankrike, men södra Frankrike var fortfarande inte fritt.
Det styrdes av "Vichy"-fransmännen. Det var fransmän som hade slutit fred med tyskarna 1940 och arbetade med inkräktarna istället för att bekämpa dem.
Den 15 augusti 1940 invaderade de allierade södra Frankrike, invasionen kallades "Operation Dragoon".
På bara två veckor hade amerikanerna och de fria franska styrkorna befriat södra Frankrike och vände sig mot Tyskland.
En civilisation är en unik kultur som delas av en betydande stor grupp människor som lever och arbetar tillsammans, ett samhälle.
Ordet civilisation kommer från latinets civilis, som betyder civil, besläktat med latinets civis, som betyder medborgare, och civitas, som betyder stad eller stadsstat, och som också på något sätt definierar samhällets storlek.
Stadsstater är föregångare till nationer. En civilisationskultur innebär att kunskap förs vidare över flera generationer, ett kvardröjande kulturellt fotavtryck och rättvis spridning.
Mindre kulturer försvinner ofta utan att lämna relevanta historiska bevis och misslyckas med att erkännas som riktiga civilisationer.
Under revolutionskriget bildade de tretton delstaterna för första gången en svag centralregering – med kongressen som enda beståndsdel – under konfederationsartiklarna.
Kongressen saknade all makt att införa skatter, och eftersom det inte fanns någon nationell verkställande eller dömande makt förlitade den sig på att statliga myndigheter, som ofta var osamarbetsvilliga, skulle genomdriva alla sina lagar.
Den hade inte heller någon befogenhet att åsidosätta skattelagar och tariffer mellan stater.
Artiklarna krävde enhälligt samtycke från alla stater innan de kunde ändras och staterna tog så lätt på centralregeringen att deras representanter ofta var frånvarande.
Italiens fotbollslandslag är tillsammans med det tyska fotbollslandslaget det näst mest framgångsrika laget i världen och blev världsmästare i fotboll 2006.
Populära sporter är fotboll, basket, volleyboll, vattenpolo, fäktning, rugby, cykling, ishockey, rullhockey och F1-motorsport.
Vintersporter är mest populära i de norra regionerna, med italienare som tävlar i internationella spel och olympiska evenemang.
Japan har nästan 7 000 öar (den största är Honshu), vilket gör Japan till den 7:e största ön i världen!
På grund av det kluster/den ögrupp som Japan har, kallas Japan ofta, på grund av sin geografiska ställning, för en "ögrupp"
Taiwan började redan på 1400-talet där europeiska sjömän som passerade förbi registrerade öns namn som Ilha Formosa, eller vacker ö.
År 1624 etablerar Nederländska Ostindiska Kompaniet en bas i sydvästra Taiwan, vilket initierar en omvandling av aboriginernas spannmålsproduktionsmetoder och anställer kinesiska arbetare för att arbeta på dess ris- och sockerplantager.
År 1683 tog Qingdynastins (1644-1912) styrkor kontroll över Taiwans västra och norra kustområden och utropade Taiwan till en provins i Qingriket 1885.
År 1895, efter nederlag i det första kinesisk-japanska kriget (1894-1895), undertecknar Qingregeringen Shimonosekifördraget, genom vilket den överlåter suveräniteten över Taiwan till Japan, som styr ön fram till 1945.
Machu Picchu består av tre huvudbyggnader, nämligen Intihuatana, Solens tempel och Rummet med de tre fönstren.
De flesta av byggnaderna i utkanten av komplexet har byggts om för att ge turisterna en bättre uppfattning om hur de ursprungligen såg ut.
År 1976 hade trettio procent av Machu Picchu restaurerats och restaureringen fortsätter än idag.
Till exempel är det vanligaste stillbildsfotograferingsformatet i världen 35 mm, som var den dominerande filmstorleken i slutet av den analoga filmeran.
Den tillverkas fortfarande idag, men ännu viktigare är att dess bildförhållande har ärvts av bildsensorformat för digitalkameror.
35 mm-formatet är faktiskt, något förvirrande, 36 mm i bredd och 24 mm i höjd.
Bildförhållandet för detta format (dividera med tolv för att få det enklaste heltalsförhållandet) sägs därför vara 3:2.
Många vanliga format (t.ex. APS-formatfamiljen) är lika med eller ligger nära det här bildförhållandet.
Den mycket missbrukade och ofta förlöjligade tredjedelsregeln är en enkel riktlinje som skapar dynamik samtidigt som den håller ett visst mått av ordning i en bild.
Den anger att den mest effektiva platsen för huvudmotivet är i skärningspunkten mellan linjer som delar bilden i tredjedelar vertikalt och horisontellt (se exempel).
Under denna period i Europas historia hamnade den katolska kyrkan, som hade blivit rik och mäktig, under lupp.
I över tusen år hade den kristna religionen bundit samman de europeiska staterna trots skillnader i språk och seder. Jag
Dess allt genomsyrande makt påverkade alla, från kung till ofrälse.
En av de viktigaste kristna grundsatserna är att rikedom ska användas för att lindra lidande och fattigdom och att kyrkans penningmedel finns där just av den anledningen.
Kyrkans centrala auktoritet hade funnits i Rom i över tusen år och denna koncentration av makt och pengar fick många att ifrågasätta om denna princip uppfylldes.
Strax efter krigsutbrottet inledde Storbritannien en sjöblockad mot Tyskland.
Strategin visade sig vara effektiv och skar av viktiga militära och civila förnödenheter, även om blockaden bröt mot allmänt accepterad internationell rätt som kodifierats av flera internationella avtal under de senaste två århundradena.
Storbritannien minerade internationellt vatten för att hindra fartyg från att komma in i hela oceaner, vilket orsakade fara även för neutrala fartyg.
Eftersom reaktionen på denna taktik var begränsad, förväntade sig Tyskland ett liknande svar på sitt obegränsade ubåtskrig.
Under 1920-talet var den förhärskande attityden hos de flesta medborgare och nationer pacifism och isolering.
Efter att ha sett krigets fasor och grymheter under första världskriget ville nationerna undvika en sådan situation igen i framtiden.
År 1884 flyttade Tesla till USA för att ta ett jobb på Edison Company i New York City.
Han anlände till USA med 4 cent i sitt namn, en poesibok och ett rekommendationsbrev från Charles Batchelor (hans manager på hans tidigare jobb) till Thomas Edison.
Det forntida Kina hade ett unikt sätt att visa olika tidsperioder; varje steg i Kina eller varje familj som satt vid makten var en distinkt dynasti.
Mellan varje dynasti rådde också en instabil tid med delade provinser. Den mest kända av dessa perioder var de tre kungadömenas epok som ägde rum i 60 år mellan Han- och Jindynastin.
Under dessa perioder utkämpades hårda strider mellan många adelsmän som stred om tronen.
De tre kungadömena var en av de blodigaste epokerna i det forntida Kinas historia, tusentals människor dog när de kämpade för att få sitta på den högsta platsen i det stora palatset i Xi'an.
Det finns många sociala och politiska effekter som användningen av metriska system, ett skifte från absolutism till republikanism, nationalism och tron på att landet tillhör folket och inte en enda härskare.
Även efter revolutionen var yrkena öppna för alla manliga sökande, vilket gjorde det möjligt för de mest ambitiösa och framgångsrika att lyckas.
Samma sak gäller för militären, för istället för att arméns rangordning baserades på klass baserades de nu på cailaber.
Den franska revolutionen inspirerade också många andra förtryckta arbetarklassmänniskor i andra länder att starta sina egna revolutioner.
Muhammed var djupt intresserad av frågor bortom detta vardagliga liv. Han brukade besöka en grotta som blev känd som "Hira" på berget "Noor" (ljus) för kontemplation.
Själva grottan, som överlevde tiderna, ger en mycket levande bild av Muhammeds andliga böjelser.
Grottan ligger på toppen av ett av bergen norr om Mecka och är helt isolerad från resten av världen.
Faktum är att det inte alls är lätt att hitta även om man visste att det fanns. Väl inne i grottan är det en total isolering.
Ingenting kan ses annat än den klara, vackra himlen ovanför och de många omgivande bergen. Väldigt lite av denna värld kan ses eller höras inifrån grottan.
Den stora pyramiden i Giza är det enda av de sju underverken som fortfarande står kvar idag.
Den stora pyramiden byggdes av egyptierna på 200-talet f.Kr. och är en av många stora pyramidstrukturer som byggdes för att hedra den döde farao.
Gizaplatån, eller "Giza-nekropolen" i den egyptiska dödsdalen innehåller flera pyramider (varav den stora pyramiden är den största), flera små gravar, flera tempel och den stora sfinxen.
Den stora pyramiden skapades för att hedra farao Khufu, och många av de mindre pyramiderna, gravarna och templen byggdes för att hedra Khufus fruar och familjemedlemmar.
"Övre bågen"-märket ser ut som ett V och "nedre bågmärket" som en häftklammer eller en fyrkant som saknar undersidan.
Upp betyder att du ska börja i spetsen och trycka på bågen, och ner betyder att du ska börja vid grodan (vilket är där din hand håller bågen) och dra bågen.
En up-bow genererar vanligtvis ett mjukare ljud, medan en down-bow är starkare och mer självsäker.
Rita gärna in dina egna märken, men kom ihåg att de tryckta stråkmärkena finns där av en musikalisk anledning, så de bör oftast respekteras.
Den skräckslagne kung Ludvig XVI, drottning Marie Antoinette, deras två små barn (11-åriga Marie Therese och fyraåriga Louis-Charles) och kungens syster, fru Elisabeth, tvingades den 6 oktober 1789 tillbaka till Paris från Versailles av en mobb av marknadskvinnor.
I en vagn färdades de tillbaka till Paris omgivna av en folkmassa som skrek och skrek hotelser mot kungen och drottningen.
Folkmassan tvingade kungen och drottningen att ha sina vagnsfönster vidöppna.
Vid ett tillfälle viftade en medlem av mobben med huvudet på en kunglig vakt som dödats i Versailles framför den skräckslagna drottningen.
USA-imperialismens krigsutgifter i samband med erövringen av Filippinerna betalades av det filippinska folket självt.
De var tvungna att betala skatt till den amerikanska kolonialregimen för att täcka en stor del av utgifterna och räntan på obligationer som flöt i den filippinska regeringens namn genom Wall Streets bankhus.
Naturligtvis skulle de superprofiter som härrör från den utdragna exploateringen av det filippinska folket utgöra de grundläggande vinsterna för USA-imperialismen.
För att förstå tempelriddarna måste man förstå det sammanhang som föranledde skapandet av orden.
Tiden då händelserna ägde rum brukar kallas högmedeltiden, den period i Europas historia under 1000-, 1100- och 1200-talen (1000–1300 e.Kr.).
Högmedeltiden föregicks av tidig medeltid och följdes av senmedeltid, som enligt konvention slutar omkring 1500.
Teknologisk determinism är en term som omfattar ett brett spektrum av idéer i praktiken, från teknik-push eller det tekniska imperativet till en strikt känsla av att människans öde drivs av en underliggande logik som är förknippad med vetenskapliga lagar och deras manifestation i teknik.
De flesta tolkningar av teknologisk determinism delar två allmänna idéer: att teknologins utveckling i sig följer en väg som till stor del går bortom kulturellt eller politiskt inflytande, och att teknologi i sin tur har "effekter" på samhällen som är medfödda, snarare än socialt betingade.
Man kan till exempel säga att bilen med nödvändighet leder till att vägar utvecklas.
Ett rikstäckande vägnät är dock inte ekonomiskt lönsamt för bara en handfull bilar, så nya produktionsmetoder utvecklas för att minska kostnaderna för bilägande.
Massägande av bilar leder också till en högre förekomst av olyckor på vägarna, vilket leder till att nya tekniker uppfinns inom sjukvården för att reparera skadade kroppar.
Romantiken hade ett stort inslag av kulturell determinism, hämtad från författare som Goethe, Fichte och Schlegel.
I samband med romantiken formade geografin individerna, och med tiden uppstod seder och bruk och kultur relaterade till denna geografi, och dessa, som var i harmoni med samhällets plats, var bättre än godtyckligt påtvingade lagar.
På samma sätt som Paris är känt som modehuvudstaden i den samtida världen, betraktades Konstantinopel som modehuvudstaden i det feodala Europa.
Dess rykte om att vara ett epicentrum för lyx började omkring 400 e.Kr. och varade fram till cirka 1100 e.Kr.
Dess status sjönk under 1100-talet, främst på grund av att korsfararna hade återvänt med gåvor som siden och kryddor som värderades högre än vad de bysantinska marknaderna erbjöd.
Det var vid denna tid som titeln modehuvudstad överfördes från Konstantinopel till Paris.
Den gotiska stilen nådde sin höjdpunkt under perioden mellan 900-1000-talet och 1300-talet.
I början var klädseln starkt influerad av den bysantinska kulturen i öst.
Men på grund av de långsamma kommunikationskanalerna kan stilar i väst släpa efter med 25 till 30 år.
Mot slutet av medeltiden började Västeuropa utveckla sin egen stil. En av de största utvecklingarna på den tiden som ett resultat av korstågen var att människor började använda knappar för att fästa kläder.
Självhushållsjordbruk är jordbruk som utförs för att producera tillräckligt med mat för att tillgodose jordbrukarens och hans/hennes familjs behov.
Självhushållande jordbruk är ett enkelt, ofta ekologiskt, system som använder sparat utsäde som är inhemskt i ekoregionen i kombination med växelbruk eller andra relativt enkla tekniker för att maximera avkastningen.
Historiskt sett har de flesta jordbrukare ägnat sig åt självhushållsjordbruk och detta är fortfarande fallet i många utvecklingsländer.
Subkulturer för samman likasinnade individer som känner sig försummade av samhällets normer och låter dem utveckla en känsla av identitet.
Subkulturer kan vara distinkta på grund av medlemmarnas ålder, etnicitet, klass, plats och/eller kön.
De kvaliteter som definierar en subkultur som distinkt kan vara språkliga, estetiska, religiösa, politiska, sexuella, geografiska eller en kombination av faktorer.
Medlemmar av en subkultur signalerar ofta sitt medlemskap genom en distinkt och symbolisk användning av stil, som inkluderar mode, manér och argot.
En av de vanligaste metoderna som används för att illustrera vikten av socialisering är att använda sig av de få olyckliga fall av barn som på grund av försummelse, olycka eller uppsåtliga övergrepp inte socialiserades av vuxna under sin uppväxt.
Sådana barn kallas "förvildade" eller vilda. En del förvildade barn har hållits instängda av människor (vanligtvis sina egna föräldrar); I vissa fall berodde övergivandet av barn på att föräldrarna avvisade ett barns allvarliga intellektuella eller fysiska funktionsnedsättning.
Förvildade barn kan ha upplevt allvarlig barnmisshandel eller trauma innan de övergavs eller rymde.
Andra påstås ha fötts upp av djur; En del sägs ha levt i det vilda på egen hand.
När det vilda barnet helt och hållet uppfostras av icke-mänskliga djur, uppvisar det beteenden (inom fysiska gränser) som nästan helt och hållet liknar det hos det särskilda djuret, såsom dess rädsla för eller likgiltighet för människor.
Även om projektbaserat lärande bör göra lärandet enklare och mer intressant, går byggnadsställningar ett steg längre.
Scaffolding är inte en metod för inlärning utan snarare ett hjälpmedel som ger stöd till individer som genomgår en ny inlärningsupplevelse som att använda ett nytt datorprogram eller påbörja ett nytt projekt.
Byggnadsställningar kan vara både virtuella och verkliga, med andra ord är en lärare en form av byggnadsställning, men det är också den lilla gemmannen i Microsoft Office.
Virtuella ställningar är internaliserade i programvaran och är avsedda att ifrågasätta, uppmana och förklara procedurer som kan ha varit för utmanande för studenten att hantera ensam.
Barn placeras i fosterhem av en mängd olika skäl som sträcker sig från försummelse, till övergrepp och till och med till utpressning.
Inget barn ska någonsin behöva växa upp i en miljö som inte är omhändertagande, omtänksam och pedagogisk, men det gör de.
Vi uppfattar familjehemssystemet som en trygghetszon för dessa barn.
Vårt fosterhemssystem är tänkt att ge trygga hem, kärleksfulla vårdgivare, stabil utbildning och pålitlig hälsovård.
Fosterhem är tänkt att tillhandahålla alla de förnödenheter som saknades i det hem de tidigare togs från.
Internet kombinerar element av både masskommunikation och interpersonell kommunikation.
Internets distinkta egenskaper leder till ytterligare dimensioner när det gäller användning och tillfredsställelse.
Till exempel föreslås "inlärning" och "socialisering" som viktiga motiv för Internetanvändning (James et al., 1995).
"Personligt engagemang" och "fortsatta relationer" identifierades också som nya motivationsaspekter av Eighmey och McCord (1998) när de undersökte publikens reaktioner på webbplatser.
Användningen av videoinspelning har lett till viktiga upptäckter i tolkningen av mikrouttryck, ansiktsrörelser som varar några millisekunder.
I synnerhet påstås det att man kan upptäcka om en person ljuger genom att tolka mikrouttryck korrekt.
Oliver Sacks visade i sin uppsats The President's Speech hur människor som inte kan förstå tal på grund av hjärnskada ändå kan bedöma uppriktighet korrekt.
Han föreslår till och med att sådana förmågor när det gäller att tolka mänskligt beteende kan delas av djur som tamhundar.
1900-talets forskning har visat att det finns två pooler av genetisk variation: dold och uttryckt.
Mutation lägger till ny genetisk variation, och selektion tar bort den från poolen av uttryckt variation.
Segregation och rekombination blandar variationen fram och tillbaka mellan de två poolerna med varje generation.
Ute på savannen är det svårt för en primat med ett matsmältningssystem som människan att tillfredsställa sitt aminosyrabehov från tillgängliga växtresurser.
Att inte göra det får dessutom allvarliga konsekvenser: tillväxtdepression, undernäring och slutligen död.
De mest lättillgängliga växtresurserna skulle ha varit de proteiner som finns i blad och baljväxter, men dessa är svåra för primater som oss att smälta om de inte är kokta.
Däremot är animaliska livsmedel (myror, termiter, ägg) inte bara lättsmälta, utan de ger också stora mängder proteiner som innehåller alla essentiella aminosyror.
Sammantaget skulle vi inte bli förvånade om våra egna förfäder löste sitt "proteinproblem" på ungefär samma sätt som schimpanserna på savannen gör idag.
Sömnavbrott är processen att målmedvetet vakna under din normala sömnperiod och somna en kort tid senare (10–60 minuter).
Detta kan enkelt göras genom att använda en relativt tyst väckarklocka för att få dig till medvetande utan att väcka dig helt.
Om du kommer på dig själv med att ställa om klockan i sömnen kan den placeras på andra sidan rummet, vilket tvingar dig att gå upp ur sängen för att stänga av den.
Andra biorytmbaserade alternativ innebär att man dricker mycket vätska (särskilt vatten eller te, ett känt diuretikum) före sömnen, vilket tvingar en att gå upp för att kissa.
Mängden inre frid som en person besitter korrelerar motsatt med mängden spänning i ens kropp och själ.
Ju lägre spänning, desto mer positiv livskraft finns. Varje person har potential att finna absolut frid och tillfredsställelse.
Alla kan uppnå upplysning. Det enda som står i vägen för detta mål är vår egen spänning och negativitet.
Den tibetanska buddhismen är baserad på Buddhas läror, men utökades av mahayana-kärlekens väg och av många tekniker från indisk yoga.
I princip är den tibetanska buddhismen mycket enkel. Den består av kundaliniyoga, meditation och den allomfattande kärlekens väg.
Med Kundaliniyoga väcks Kundalinienergin (upplysningsenergin) genom yogaställningar, andningsövningar, mantran och visualiseringar.
Centrum för tibetansk meditation är gudomsyogan. Genom visualisering av olika gudar renas energikanalerna, chakrana aktiveras och upplysningsmedvetandet skapas.
Tyskland var en gemensam fiende i andra världskriget, vilket ledde till samarbete mellan Sovjetunionen och USA. I och med krigsslutet ledde konflikterna mellan system, processer och kultur till att länderna föll osams.
Med två år efter krigsslutet var de tidigare allierade nu fiender och det kalla kriget började.
Den skulle pågå under de kommande 40 åren och skulle utkämpas på riktigt, av proxyarméer, på slagfält från Afrika till Asien, i Afghanistan, Kuba och på många andra platser.
Den 17 september 1939 var det polska försvaret redan brutet, och det enda hoppet var att dra sig tillbaka och omorganisera sig längs det rumänska brohuvudet.
Dessa planer blev dock föråldrade nästan över en natt, när över 800 000 soldater från Sovjetunionens Röda armé gick in och skapade de vitryska och ukrainska fronterna efter att ha invaderat de östra regionerna i Polen i strid med fredsfördraget i Riga, den sovjetisk-polska icke-angreppspakten och andra internationella fördrag, både bilaterala och multilaterala.
Att använda fartyg för att transportera varor är det överlägset mest effektiva sättet att flytta stora mängder människor och varor över haven.
Flottornas uppgift har traditionellt varit att se till att ditt land behåller förmågan att flytta ditt folk och dina varor, samtidigt som du stör din fiendes förmåga att flytta sitt folk och sina varor.
Ett av de mest anmärkningsvärda exemplen på detta på senare tid var den nordatlantiska kampanjen under andra världskriget. Amerikanerna försökte transportera män och material över Atlanten för att hjälpa Storbritannien.
Samtidigt försökte den tyska flottan, främst med hjälp av ubåtar, stoppa denna trafik.
Om de allierade hade misslyckats skulle Tyskland förmodligen ha kunnat erövra Storbritannien på samma sätt som resten av Europa.
Getter verkar ha domesticerats för ungefär 10 000 år sedan i Zagrosbergen i Iran.
Forntida kulturer och stammar började hålla dem för att de skulle vara lätta att få tillgång till mjölk, hår, kött och skinn.
Tamgetter hölls i allmänhet i hjordar som vandrade på kullar eller andra betesmarker, ofta skötta av getherdar som ofta var barn eller ungdomar, liknande den mer allmänt kända herden. Dessa metoder används än idag.
Vagnvägar byggdes i England redan på 1500-talet.
Även om vagnbanorna bara bestod av parallella träplankor, tillät de hästar som drog dem att uppnå högre hastigheter och dra större laster än på de lite mer ojämna vägarna på den tiden.
Korsband infördes ganska tidigt för att hålla spåren på plats. Så småningom insåg man dock att banden skulle bli mer effektiva om de hade en järnspets på toppen.
Detta blev vanligt förekommande, men järnet orsakade mer slitage på vagnarnas trähjul.
Så småningom ersattes trähjul av järnhjul. År 1767 introducerades de första rälsen av heljärn.
Den första kända transporten var att gå, människor började gå upprätt för två miljoner år sedan med uppkomsten av Homo Erectus (som betyder upprätt människa).
Deras föregångare, Australopithecus, gick inte upprätt som vanligt.
Tvåbenta specialiseringar har hittats i fossil av Australopithecus för 4,2-3,9 miljoner år sedan, även om Sahelanthropus kan ha gått på två ben så tidigt som för sju miljoner år sedan.
Vi kan börja leva mer miljövänligt, vi kan gå med i miljörörelsen och vi kan till och med vara aktivister för att minska det framtida lidandet i viss mån.
Detta är i många fall precis som symtomatisk behandling. Men om vi inte bara vill ha en tillfällig lösning bör vi hitta roten till problemen, och vi bör inaktivera dem.
Det är uppenbart nog att världen har förändrats mycket på grund av mänsklighetens vetenskapliga och tekniska framsteg, och problemen har blivit större på grund av överbefolkning och mänsklighetens extravaganta livsstil.
Efter att det antagits av kongressen den 4 juli skickades ett handskrivet utkast undertecknat av kongressens ordförande John Hancock och sekreteraren Charles Thomson några kvarter bort till John Dunlaps tryckeri.
Under natten tillverkades mellan 150 och 200 exemplar, numera kända som "Dunlap broadsides".
Den första offentliga uppläsningen av dokumentet gjordes av John Nixon på gården till Independence Hall den 8 juli.
En sändes till George Washington den 6 juli, som fick den uppläst för sina trupper i New York den 9 juli. En kopia nådde London den 10 augusti.
De 25 Dunlap-skillingtryck som fortfarande finns kvar är de äldsta bevarade kopiorna av dokumentet. Den handskrivna originalkopian har inte överlevt.
Många paleontologer tror idag att en grupp dinosaurier överlevde och lever idag. Vi kallar dem fåglar.
Många tänker inte på dem som dinosaurier eftersom de har fjädrar och kan flyga.
Men det finns många saker med fåglar som fortfarande ser ut som en dinosaurie.
De har fötter med fjäll och klor, de lägger ägg och de går på sina två bakben som en T-Rex.
I stort sett alla datorer som används idag bygger på manipulation av information som är kodad i form av binära tal.
Ett binärt tal kan bara ha ett av två värden, dvs. 0 eller 1, och dessa tal kallas binära siffror - eller bitar, för att använda datorjargong.
Inre förgiftning kanske inte är omedelbart uppenbar. Symtomen, såsom kräkningar, är tillräckligt allmänna för att en omedelbar diagnos inte ska kunna ställas.
Den bästa indikationen på intern förgiftning kan vara närvaron av en öppen behållare med läkemedel eller giftiga hushållskemikalier.
Kontrollera etiketten för specifika första hjälpen-instruktioner för det specifika giftet.
Termen insekt används av entomologer i formell bemärkelse för denna grupp av insekter.
Denna term härstammar från forntida förtrogenhet med vägglöss, som är insekter som är mycket anpassade för att parasitera människor.
Både lönnmördarbaggar och vägglöss är nidicolous, anpassade till att leva i bo eller bostad hos sin värd.
I USA finns det cirka 400 000 kända fall av multipel skleros (MS), vilket gör den till den ledande neurologiska sjukdomen hos yngre och medelålders vuxna.
MS är en sjukdom som påverkar det centrala nervsystemet, som består av hjärnan, ryggmärgen och synnerven.
Forskning har visat att kvinnor löper två gånger större risk att få MS än män.
Ett par kan bestämma sig för att det inte är i deras eget intresse, eller i deras barns intresse, att uppfostra ett barn.
Dessa par kan välja att göra en adoptionsplan för sitt barn.
Vid en adoption upphäver de biologiska föräldrarna sina föräldrarättigheter så att ett annat par kan ta hand om barnet.
Vetenskapens huvudmål är att ta reda på hur världen fungerar genom den vetenskapliga metoden. Denna metod vägleder i själva verket den mesta vetenskapliga forskningen.
Det är dock inte ensamt, experiment, och ett experiment är ett test som används för att eliminera en eller flera av de möjliga hypoteserna, ställa frågor och göra observationer vägleder också vetenskaplig forskning.
Naturforskare och filosofer fokuserade på klassiska texter och i synnerhet på Bibeln på latin.
Aristoteles åsikter om alla vetenskapliga frågor, inklusive psykologi, accepterades.
I takt med att kunskaperna i grekiska minskade, fann sig västvärlden avskuren från sina grekiska filosofiska och vetenskapliga rötter.
Många observerade rytmer i fysiologi och beteende beror ofta på närvaron av endogena cykler och deras produktion genom biologiska klockor.
Periodiska rytmer, som inte bara är svar på externa periodiska signaler, har dokumenterats för de flesta levande varelser, inklusive bakterier, svampar, växter och djur.
Biologiska klockor är självförsörjande oscillatorer som kommer att fortsätta en period av fritt springande cykling även i frånvaro av externa signaler.
Hershey och Chase-experimentet var ett av de ledande förslagen om att DNA var ett genetiskt material.
Hershey och Chase använde fager, eller virus, för att implantera sitt eget DNA i en bakterie.
De gjorde två experiment där de antingen markerade DNA i fagen med en radioaktiv fosfor eller fagens protein med radioaktivt svavel.
Mutationer kan ha en mängd olika effekter beroende på vilken typ av mutation det rör sig om, vilken betydelse det genetiska materialet har och om de celler som påverkas är könsceller.
Endast mutationer i könsceller kan föras vidare till barn, medan mutationer på andra håll kan orsaka celldöd eller cancer.
Naturbaserad turism lockar människor som är intresserade av att besöka naturområden i syfte att njuta av landskapet, inklusive växt- och djurliv.
Exempel på aktiviteter på plats är jakt, fiske, fotografering, fågelskådning och besök i parker och studier av information om ekosystemet.
Ett exempel är att besöka, fotografera och lära sig om organgatuangs på Borneo.
Varje morgon lämnar människor små landsortsstäder i bilar för att åka till sin arbetsplats och blir omkörda av andra vars arbetsplats är den plats de just har lämnat.
I denna dynamiska transportbuss är alla på något sätt anslutna till och stöder ett transportsystem baserat på privatbilar.
Vetenskapen visar nu att denna massiva kolekonomi har förskjutit biosfären från ett av dess stabila tillstånd som har stött människans evolution under de senaste två miljoner åren.
Alla deltar i samhället och använder transportsystem. Nästan alla klagar på transportsystemen.
I utvecklade länder hör man sällan liknande nivåer av klagomål om vattenkvalitet eller broar som rasar.
Varför ger transportsystemen upphov till sådana klagomål, varför misslyckas de dagligen? Är transportingenjörer bara inkompetenta? Eller är det något mer grundläggande som pågår?
Trafikflöde är studiet av enskilda förares och fordons rörelse mellan två punkter och de interaktioner de gör med varandra.
Tyvärr är det svårt att studera trafikflödet eftersom förarens beteende inte kan förutsägas med hundra procents säkerhet.
Lyckligtvis tenderar förare att bete sig inom ett någorlunda konsekvent intervall; Trafikströmmar tenderar därför att ha en rimlig konsekvens och kan grovt representeras matematiskt.
För att bättre representera trafikflödet har samband etablerats mellan de tre huvudegenskaperna: (1) flöde, (2) densitet och (3) hastighet.
Dessa relationer hjälper till vid planering, design och drift av väganläggningar.
Insekter var de första djuren som tog sig upp i luften. Deras förmåga att flyga hjälpte dem att lättare undvika fiender och hitta mat och partners mer effektivt.
De flesta insekter har fördelen att kunna fälla tillbaka vingarna längs kroppen.
Detta ger dem ett större utbud av små platser att gömma sig från rovdjur.
Idag är de enda insekter som inte kan fälla tillbaka sina vingar trollsländor och dagsländor.
För tusentals år sedan sa en man vid namn Aristarchos att solsystemet rörde sig runt solen.
En del trodde att han hade rätt, men många trodde motsatsen. att solsystemet rörde sig runt jorden, inklusive solen (och till och med de andra stjärnorna).
Detta verkar vettigt, för det känns inte som om jorden rör sig, eller hur?
Amazonfloden är den näst längsta och största floden på jorden. Den bär mer än 8 gånger så mycket vatten som den näst största floden.
Amazonas är också den bredaste floden på jorden, ibland sex mil bred.
Hela 20 procent av det vatten som rinner ut ur planetens floder i haven kommer från Amazonas.
Amazonflodens huvudflod är 6 387 km (3 980 miles). Den samlar upp vatten från tusentals mindre floder.
Även om pyramidbyggandet i sten fortsatte fram till slutet av Gamla riket, överträffades pyramiderna i Giza aldrig i sin storlek och den tekniska förträffligheten i deras konstruktion.
Nya rikets forntida egyptier förundrades över sina föregångares monument, som då var långt över tusen år gamla.
Vatikanstaten har cirka 800 invånare. Det är det minsta självständiga landet i världen och det land som har lägst befolkning.
Vatikanstaten använder italienska i sin lagstiftning och officiella kommunikation.
Italienska är också det vardagsspråk som används av de flesta som arbetar i staten, medan latin ofta används i religiösa ceremonier.
Alla medborgare i Vatikanstaten är romersk-katolska.
Människor har känt till grundläggande kemiska grundämnen som guld, silver och koppar sedan antiken, eftersom dessa alla kan upptäckas i naturen i inhemsk form och är relativt enkla att bryta med primitiva verktyg.
Aristoteles, en filosof, teoretiserade att allt består av en blandning av ett eller flera av fyra element. De var jord, vatten, luft och eld.
Detta var mer likt de fyra materiens tillstånd (i samma ordning): fast, flytande, gas och plasma, även om han också teoretiserade att de förändras till nya ämnen för att bilda det vi ser.
Legeringar är i grunden en blandning av två eller flera metaller. Glöm inte att det finns många grundämnen i det periodiska systemet.
Grundämnen som kalcium och kalium anses vara metaller. Naturligtvis finns det också metaller som silver och guld.
Du kan också ha legeringar som innehåller små mängder icke-metalliska element som kol.
Allting i universum är gjort av materia. All materia består av små partiklar som kallas atomer.
Atomer är så otroligt små att biljoner av dem skulle kunna passa in i perioden i slutet av den här meningen.
Pennan var alltså en god vän till många människor när den kom ut.
Tyvärr, i takt med att nyare skrivmetoder har dykt upp, har pennan förpassats till mindre status och användningsområden.
Människor skriver nu meddelanden på datorskärmar och behöver aldrig komma i närheten av en vässare.
Man kan bara undra vad tangentbordet kommer att bli när något nyare dyker upp.
Fissionsbomben fungerar enligt principen att det krävs energi för att sätta ihop en kärna med många protoner och neutroner.
Ungefär som att rulla en tung vagn uppför en backe. Att dela upp kärnan igen frigör då en del av den energin.
Vissa atomer har instabila kärnor vilket innebär att de tenderar att brytas isär med liten eller ingen knuff.
Månens yta är gjord av stenar och stoft. Månens yttre lager kallas skorpan.
Jordskorpan är ca 70 km tjock på den närmaste sidan och 100 km tjock på den bortre sidan.
Den är tunnare under marian och tjockare under höglandet.
Det kan finnas mer maria på den närmaste sidan eftersom skorpan är tunnare. Det var lättare för lava att stiga upp till ytan.
Innehållsteorier är inriktade på att hitta det som får människor att ticka eller tilltalar dem.
Dessa teorier föreslår att människor har vissa behov och/eller önskningar som har internaliserats när de mognar till vuxen ålder.
Dessa teorier tittar på vad det är med vissa personer som får dem att vilja ha de saker de gör och vilka saker i deras omgivning som får dem att göra eller inte göra vissa saker.
Två populära innehållsteorier är Maslows behovshierarkiteori och Hertzbergs tvåfaktorteori.
Generellt sett kan två beteenden uppstå när chefer börjar leda sina tidigare kollegor. Ena änden av spektrumet är att försöka förbli "en av killarna" (eller tjejerna).
Denna typ av chef har svårt att fatta impopulära beslut, utföra disciplinära åtgärder, prestationsutvärderingar, tilldela ansvar och hålla människor ansvariga.
I andra änden av spektrumet förvandlas en till en oigenkännlig individ som känner att han eller hon måste ändra allt som teamet har gjort och göra det till sitt eget.
När allt kommer omkring är ledaren ytterst ansvarig för teamets framgång och misslyckande.
Detta beteende resulterar ofta i sprickor mellan ledarna och resten av teamet.
Virtuella team håller samma standarder för excellens som konventionella team, men det finns subtila skillnader.
Virtuella teammedlemmar fungerar ofta som kontaktpunkt för sin närmaste fysiska grupp.
De har ofta mer självständighet än konventionella teammedlemmar eftersom deras team kan träffas enligt olika tidszoner som kanske inte förstås av deras lokala ledning.
Närvaron av ett verkligt "osynligt team" (Larson och LaFasto, 1989, s109) är också en unik komponent i ett virtuellt team.
Det "osynliga teamet" är den ledningsgrupp som var och en av medlemmarna rapporterar till. Det osynliga teamet sätter standarden för varje medlem.
Varför skulle en organisation vilja gå igenom den tidskrävande processen att etablera en lärande organisation? Ett mål för att omsätta organisatoriska inlärningskoncept i praktiken är innovation.
När alla tillgängliga resurser används effektivt på de funktionella avdelningarna i en organisation kan kreativitet och uppfinningsrikedom uppstå.
Som ett resultat kan processen för en organisation som arbetar tillsammans för att övervinna ett hinder leda till en ny innovativ process för att tillgodose kundens behov.
Innan en organisation kan vara innovativ måste ledarskapet skapa en kultur av innovation samt delad kunskap och organisatoriskt lärande.
Angel (2006) förklarar Continuum-metoden som en metod som används för att hjälpa organisationer att nå en högre prestationsnivå.
Neurobiologiska data ger fysiska bevis för ett teoretiskt tillvägagångssätt för att undersöka kognition. Därför begränsar det forskningsområdet och gör det mycket mer exakt.
Sambandet mellan hjärnpatologi och beteende stöder forskare i deras forskning.
Det har länge varit känt att olika typer av hjärnskador, trauman, skador och tumörer påverkar beteendet och orsakar förändringar i vissa mentala funktioner.
Framväxten av ny teknik gör det möjligt för oss att se och undersöka hjärnstrukturer och processer som aldrig tidigare skådats.
Detta ger oss mycket information och material för att bygga simuleringsmodeller som hjälper oss att förstå processer i vårt sinne.
Även om AI har en stark koppling till science fiction utgör AI en mycket viktig gren av datavetenskapen, som handlar om beteende, inlärning och intelligent anpassning i en maskin.
Forskning inom AI handlar om att få maskiner att automatisera uppgifter som kräver intelligent beteende.
Exempel på detta är kontroll, planering och schemaläggning, förmågan att svara på kunddiagnoser och frågor samt handskriftsigenkänning, röst och ansikte.
Sådana saker har blivit separata discipliner, som fokuserar på att tillhandahålla lösningar på verkliga problem.
AI-systemet används nu ofta inom ekonomi, medicin, teknik och militär, vilket har byggts in i flera hemdator- och videospelsprogram.
Studiebesök är en stor del av alla klassrum. Ganska ofta skulle en lärare älska att ta med sina elever till platser dit en bussresa inte är ett alternativ.
Tekniken erbjuder lösningen med virtuella studiebesök. Eleverna kan titta på museiföremål, besöka ett akvarium eller beundra vacker konst medan de sitter med sin klass.
Att dela en studieresa virtuellt är också ett bra sätt att reflektera över en resa och dela erfarenheter med framtida klasser.
Till exempel designar elever från Bennet School i North Carolina varje år en webbplats om sin resa till delstatshuvudstaden, varje år görs webbplatsen om, men gamla versioner sparas online för att fungera som en klippbok.
Bloggar kan också bidra till att förbättra elevernas skrivande. Även om studenter ofta börjar sin bloggupplevelse med slarvig grammatik och stavning, ändrar närvaron av en publik i allmänhet det.
Eftersom studenter ofta är den mest kritiska publiken börjar bloggskribenten sträva efter att förbättra skrivandet för att undvika kritik.
Att blogga "tvingar också eleverna att bli mer kunniga om världen omkring dem." Behovet av att väcka publikens intresse inspirerar eleverna att vara smarta och intressanta (Toto, 2004).
Att blogga är ett verktyg som inspirerar till samarbete och uppmuntrar eleverna att utöka lärandet långt bortom den traditionella skoldagen.
Lämplig användning av bloggar "kan ge eleverna möjlighet att bli mer analytiska och kritiska; Genom att aktivt reagera på Internetmaterial kan eleverna definiera sina ståndpunkter i samband med andras skrifter samt skissera sina egna perspektiv på särskilda frågor (Oravec, 2002).
Ottawa är Kanadas charmiga, tvåspråkiga huvudstad och har en rad konstgallerier och museer som visar upp Kanadas förflutna och nutid.
Längre söderut ligger Niagarafallen och i norr finns den outnyttjade naturliga skönheten i Muskoka och bortom.
Alla dessa saker och mer därtill framhäver Ontario som vad som anses vara typiskt kanadensiskt av utomstående.
Stora områden längre norrut är ganska glesbefolkade och en del är nästan obebodd vildmark.
För en jämförelse av befolkningen som förvånar många: Det bor fler afroamerikaner i USA än det finns kanadensiska medborgare.
De östafrikanska öarna ligger i Indiska oceanen utanför Afrikas östkust.
Madagaskar är den överlägset största, och en egen kontinent när det kommer till djurliv.
De flesta av de mindre öarna är självständiga nationer, eller associerade med Frankrike, och kända som lyxiga badorter.
Araberna förde också med sig islam till länderna, och det tog stor plats på Komorerna och Mayotte.
Det europeiska inflytandet och kolonialismen började på 1400-talet, när den portugisiske upptäcktsresanden Vasco da Gama hittade Kapvägen från Europa till Indien.
I norr avgränsas regionen av Sahel och i söder och väster av Atlanten.
Kvinnor: Det rekommenderas att alla kvinnliga resenärer uppger att de är gifta, oavsett faktiskt civilstånd.
Det är bra att också bära en ring (bara inte en som ser för dyr ut.
Kvinnor bör inse att kulturella skillnader kan resultera i vad de skulle betrakta som trakasserier och det är inte ovanligt att bli förföljd, gripen i armen etc.
Var bestämd när du tackar nej till män, och var inte rädd för att stå på dig (kulturella skillnader eller inte, det gör det inte ok!).
Den moderna staden Casablanca grundades av berbiska fiskare på 900-talet f.Kr. och användes av fenicierna, romarna och mereniderna som en strategisk hamn vid namn Anfa.
Portugiserna förstörde den och återuppbyggde den under namnet Casa Branca, bara för att överge den efter en jordbävning 1755.
Den marockanska sultanen byggde om staden till Daru l-Badya och den fick namnet Casablanca av spanska handelsmän som etablerade handelsbaser där.
Casablanca är en av de minst intressanta platserna att shoppa på i hela Marocko.
Runt den gamla medinan är det lätt att hitta ställen som säljer traditionella marockanska varor, såsom tagines, keramik, lädervaror, vattenpipor och ett helt spektrum av geegaws, men allt är för turisterna.
Goma är en turiststad i Demokratiska republiken Kongo i Yttersta östern nära Rwanda.
År 2002 förstördes Goma av lava från vulkanen Nyiragongo som begravde de flesta av stadens gator, särskilt stadens centrum.
Även om Goma är någorlunda säkert, bör alla besök utanför Goma undersökas för att förstå tillståndet i striderna som fortsätter i Nordkivu-provinsen.
Staden är också basen för att bestiga vulkanen Nyiragongo tillsammans med några av de billigaste bergsgorillaspårningarna i Afrika.
Du kan använda boda-boda (motorcykeltaxi) för att ta dig runt i Goma. Det normala (lokala) priset är ~500 kongolesiska franc för den korta resan.
I kombination med sin relativa otillgänglighet har "Timbuktu" kommit att användas som en metafor för exotiska, fjärran länder.
Idag är Timbuktu en fattig stad, även om dess rykte gör den till en turistattraktion, och den har en flygplats.
År 1990 lades den till på listan över världsarv i fara på grund av hotet från ökensand.
Det var ett av de stora stoppen under Henry Louis Gates PBS-special Wonders of the African World.
Staden står i skarp kontrast till resten av landets städer, eftersom den har mer av en arabisk stil än en afrikansk.
Kruger National Park (KNP) ligger i nordöstra Sydafrika och sträcker sig längs gränsen till Moçambique i öster, Zimbabwe i norr och den södra gränsen är Crocodile River.
Parken täcker 19 500 km² och är uppdelad i 14 olika ekozoner, som var och en stöder olika vilda djur.
Det är en av Sydafrikas huvudattraktioner och anses vara flaggskeppet för sydafrikanska nationalparker (SANParks).
Som med alla sydafrikanska nationalparker finns det dagliga bevarande- och inträdesavgifter för parken.
Det kan också vara fördelaktigt för en att köpa ett Wild Card, som ger inträde till antingen urval av parker i Sydafrika eller alla de sydafrikanska nationalparkerna.
Hongkongön ger territoriet Hongkong sitt namn och är den plats som många turister betraktar som huvudfokus.
Paraden av byggnader som utgör Hongkongs skyline har liknats vid ett glittrande stapeldiagram som blir uppenbart av närvaron av vattnet i Victoria Harbour.
För att få den bästa utsikten över Hongkong, lämna ön och bege dig till Kowloons strandpromenad mittemot.
Den stora majoriteten av Hongkongöns stadsutveckling är tätt packad på återvunnen mark längs den norra kusten.
Detta är den plats som de brittiska kolonisatörerna tog som sin egen, så om du letar efter bevis på territoriets koloniala förflutna är detta ett bra ställe att börja.
Sundarbans är det största mangrovebältet i världen och sträcker sig 80 km in i Bangladeshs och Indiens inland från kusten.
Sundarbans har förklarats som ett av UNESCO:s världsarv. Den del av skogen som ligger på indiskt territorium kallas Sundarbans nationalpark.
Skogarna är dock inte bara mangroveträsk - de inkluderar några av de sista kvarvarande bestånden av de mäktiga djunglerna som en gång täckte Gangeslätten.
Sundarbans täcker en yta på 3 850 km², varav ungefär en tredjedel är täckt av vatten/träskområden.
Sedan 1966 har Sundarbans varit ett viltreservat, och det uppskattas att det nu finns 400 kungliga bengaliska tigrar och cirka 30 000 fläckiga hjortar i området.
Bussarna avgår från busstationen mellan distrikten (på andra sidan floden) under hela dagen, men de flesta, särskilt de som går österut och Jakar/Bumthang, avgår mellan 06:30 och 07:30.
Eftersom bussarna mellan distrikten ofta är fulla är det lämpligt att köpa en biljett några dagar i förväg.
De flesta distrikt betjänas av små japanska berg- och dalbanebussar, som är bekväma och robusta.
Delade taxibilar är ett snabbt och bekvämt sätt att resa till närliggande platser, till exempel Paro (Nu 150) och Punakha (Nu 200).
Oyapock River Bridge är en snedkabelbro. Den sträcker sig över floden Oyapock för att förbinda städerna Oiapoque i Brasilien och Saint-Georges de l'Oyapock i Franska Guyana.
De två tornen reser sig till en höjd av 83 meter, det är 378 meter långt och det har två filer på 3,50 m breda.
Den fria höjden under bron är 15 meter. Bygget slutfördes i augusti 2011 och öppnades inte för trafik förrän i mars 2017.
Bron är planerad att vara i full drift i september 2017, då de brasilianska tullkontrollerna förväntas vara klara.
Guaraní var den mest betydande inhemska gruppen som bodde i det som nu är östra Paraguay, och levde som halvnomadiska jägare som också utövade självhushållande jordbruk.
Chaco-regionen var hem för andra grupper av inhemska stammar som Guaycurú och Payaguá, som överlevde genom att jaga, samla och fiska.
På 1500-talet föddes Paraguay, tidigare kallat "Indiens jätteprovins", som ett resultat av de spanska erövrarnas möte med de inhemska folkgrupperna.
Spanjorerna inledde kolonisationsperioden som varade i tre århundraden.
Sedan grundandet av Asunción 1537 har Paraguay lyckats behålla mycket av sin inhemska karaktär och identitet.
Argentina är känt för att ha ett av de bästa pololagen och spelarna i världen.
Årets största turnering äger rum i december på poloplanerna i Las Cañitas.
Mindre turneringar och matcher kan även ses här under andra tider på året.
För nyheter om turneringar och var du kan köpa biljetter till polomatcher, kolla in Asociacion Argentina de Polo.
Den officiella valutan för Falklandsöarna är Falklandspund (FKP) vars värde motsvarar ett brittiskt pund (GBP).
Pengar kan växlas på den enda banken på öarna som ligger i Stanley mittemot FIC West-butiken.
Brittiska pund accepteras i allmänhet var som helst på öarna och inom Stanley accepteras ofta kreditkort och amerikanska dollar.
På de avlägsna öarna kommer kreditkort förmodligen inte att accepteras, även om brittisk och amerikansk valuta kan tas. Kontrollera med ägarna i förväg för att avgöra vad som är en acceptabel betalningsmetod.
Det är nästan omöjligt att växla Falklandsvaluta utanför öarna, så växla pengar innan du lämnar öarna.
Eftersom Montevideo ligger söder om ekvatorn är det sommar där när det är vinter på norra halvklotet och vice versa.
Montevideo ligger i subtropikerna; Under sommarmånaderna är temperaturer över +30°C vanliga.
Vintern kan vara bedrägligt kylig: temperaturen går sällan under fryspunkten, men vinden och luftfuktigheten gör att det känns kallare än vad termometern visar.
Det finns inga särskilda "regniga" och "torra" årstider: mängden regn förblir ungefär densamma under hela året.
Även om många av djuren i parken är vana vid att se människor, är djurlivet ändå vilt och bör inte matas eller störas.
Enligt parkmyndigheterna, håll dig minst 100 meter/meter från björnar och vargar och 25 meter/meter från alla andra vilda djur!
Oavsett hur fogliga de ser ut kan bisonoxar, älgar, älgar, björnar och nästan alla stora djur attackera.
Varje år skadas dussintals besökare för att de inte hållit ordentligt avstånd. Dessa djur är stora, vilda och potentiellt farliga, så ge dem deras utrymme.
Var dessutom medveten om att lukter lockar till sig björnar och andra vilda djur, så undvik att bära eller laga luktande mat och håll ett rent läger.
Apia är Samoas huvudstad. Staden ligger på ön Upolu och har en befolkning på knappt 40 000.
Apia grundades på 1850-talet och har varit Samoas officiella huvudstad sedan 1959.
Hamnen var platsen för ett ökänt sjöstillestånd 1889 när sju fartyg från Tyskland, USA och Storbritannien vägrade att lämna hamnen.
Alla fartyg sänktes, utom en brittisk kryssare. Nästan 200 amerikaner och tyskar miste livet.
Under kampen för självständighet som organiserades av Mau-rörelsen resulterade en fredlig sammankomst i staden i att den högste ledaren Tupua Tamasese Lealofi III dödades.
Det finns många stränder på grund av Aucklands gränsdragning mellan två hamnar. De mest populära finns inom tre områden.
North Shore-stränderna (i North Harbour-distriktet) ligger vid Stilla havet och sträcker sig från Long Bay i norr till Devonport i söder.
De är nästan alla sandstränder med säker simning, och de flesta har skugga från pohutukawa-träd.
Stränderna på Tamaki Drive ligger i Waitemata Harbour, i de exklusiva förorterna Mission Bay och St Heliers i centrala Auckland.
Dessa är ibland trånga familjestränder med ett bra utbud av butiker som kantar stranden. Simning är säkert.
Den viktigaste lokala ölen är "Number One", det är inte en komplex öl, men trevlig och uppfriskande. Den andra lokala ölen heter "Manta".
Det finns många franska viner att få, men de nyzeeländska och australiensiska vinerna kanske reser bättre.
Det lokala kranvattnet är helt säkert att dricka, men vatten på flaska är lätt att hitta om du är rädd.
För australiensare är tanken på "flat white" kaffe främmande. En kort svart är "espresso", cappuccino kommer hög med grädde (inte skum) och te serveras utan mjölk.
Den varma chokladen är upp till belgisk standard. Fruktjuicer är dyra men utmärkta.
Många resor till revet görs året runt, och skador på grund av någon av dessa orsaker på revet är sällsynta.
Ta ändå råd från myndigheter, följ alla skyltar och var uppmärksam på säkerhetsvarningar.
Kubmaneter förekommer nära stränder och nära flodmynningar från oktober till april norr om 1770. De kan ibland hittas utanför dessa tider.
Hajar finns, men de attackerar sällan människor. De flesta hajar är rädda för människor och skulle simma iväg.
Saltvattenkrokodiler lever inte aktivt i havet, deras primära livsmiljö är i flodmynningar norr om Rockhampton.
Att boka i förväg ger resenären sinnesfrid att de kommer att ha någonstans att sova när de anländer till sin destination.
Resebyråer har ofta avtal med specifika hotell, även om du kan tycka att det är möjligt att boka andra former av boende, som campingplatser, via en resebyrå.
Resebyråer erbjuder vanligtvis paket som inkluderar frukost, transportarrangemang till/från flygplatsen eller till och med kombinerade flyg- och hotellpaket.
De kan också hålla bokningen åt dig om du behöver tid att tänka på erbjudandet eller skaffa andra dokument för din destination (t.ex. visum).
Eventuella ändringar eller önskemål bör dock framföras via resebyrån först och inte direkt med hotellet.
För vissa festivaler bestämmer sig den stora majoriteten av deltagarna på musikfestivaler för att campa på plats, och de flesta deltagare anser att det är en viktig del av upplevelsen.
Om du vill vara nära händelsernas centrum måste du komma in tidigt för att få en campingplats nära musiken.
Kom ihåg att även om musiken på huvudscenerna kan ha slutat, kan det finnas delar av festivalen som fortsätter att spela musik till sent in på natten.
Vissa festivaler har särskilda campingområden för familjer med små barn.
Om du korsar norra Östersjön på vintern, kontrollera stugans läge, eftersom isen orsakar ganska hemskt buller för dem som drabbas hårdast.
Sankt Petersburg kryssningar inkluderar tid i stan. Kryssningspassagerare är undantagna från visumkrav (kontrollera villkoren).
Casinon gör vanligtvis många ansträngningar för att maximera den tid och de pengar som gästerna spenderar. Fönster och klockor saknas vanligtvis och utgångar kan vara svåra att hitta.
De har vanligtvis speciella mat-, dryckes- och underhållningserbjudanden för att hålla gästerna på gott humör och hålla dem i lokalen.
Vissa ställen erbjuder alkoholhaltiga drycker i huset. Fylleri försämrar dock omdömet, och alla bra spelare vet vikten av att hålla sig nykter.
Alla som ska köra på höga breddgrader eller över bergspass bör överväga möjligheten till snö, is eller minusgrader.
På isiga och snöiga vägar är friktionen låg och du kan inte köra som om du befann dig på bar asfalt.
Under snöstormar kan tillräckligt med snö falla på mycket kort tid.
Sikten kan också begränsas av fallande eller blåsande snö eller av kondens eller is på fordonsrutorna.
Å andra sidan är isiga och snöiga förhållanden normala i många länder, och trafiken pågår i stort sett oavbrutet året runt.
Safaris är kanske den största turistattraktionen i Afrika och höjdpunkten för många besökare.
Termen safari i populärt bruk hänvisar till landresor för att se det fantastiska afrikanska djurlivet, särskilt på savannen.
Vissa djur, som elefanter och giraffer, tenderar att närma sig bilar och standardutrustning gör det möjligt att se dem bra.
Lejon, geparder och leoparder är ibland skygga och du ser dem bättre med kikare.
En vandringssafari (även kallad "bush walk", "vandringssafari" eller att gå "fot") består av vandring, antingen i några timmar eller flera dagar.
Paralympics kommer att äga rum från den 24 augusti till den 5 september 2021. Vissa evenemang kommer att hållas på andra platser i Japan.
Tokyo kommer att vara den enda asiatiska staden som har varit värd för två sommar-OS, efter att ha varit värd för spelen 1964.
Om du bokade flyg och boende för 2020 innan uppskjutningen tillkännagavs kan du ha en knepig situation.
Avbokningsreglerna varierar, men från och med slutet av mars gäller de flesta avbokningsregler på grund av coronaviruset inte till juli 2020, då OS hade planerats.
Det förväntas att de flesta evenemangsbiljetter kommer att kosta mellan 2 500 och 130 000 yen, med typiska biljetter som kostar cirka 7 000 yen.
Att stryka fuktiga kläder kan hjälpa dem att torka. Många hotell har strykjärn och strykbräda att låna, även om det inte finns någon på rummet.
Om ett strykjärn inte finns tillgängligt, eller om du inte vill bära strukna strumpor, kan du prova att använda en hårtork, om tillgänglig.
Var noga med att inte låta tyget bli för varmt (vilket kan orsaka krympning eller i extrema fall sveda).
Det finns olika sätt att rena vatten, vissa mer effektiva mot specifika hot.
I vissa områden räcker det med att koka vatten i en minut, i andra behövs flera minuter.
Filter varierar i effektivitet, och om du är orolig bör du överväga att köpa ditt vatten i en förseglad flaska från ett välrenommerat företag.
Resenärer kan stöta på skadedjur som de inte känner till i sina hemtrakter.
Skadedjur kan förstöra mat, orsaka irritation eller i värsta fall orsaka allergiska reaktioner, sprida gift eller överföra infektioner.
Infektionssjukdomar i sig, eller farliga djur som kan skada eller döda människor med våld, räknas vanligtvis inte som skadedjur.
Taxfree-shopping är möjligheten att köpa varor som är befriade från skatter och punktskatter på vissa platser.
Resenärer som är på väg till länder med hög beskattning kan ibland spara en ansenlig summa pengar, särskilt på produkter som alkoholhaltiga drycker och tobak.
Sträckan mellan Point Marion och Fairmont erbjuder de mest utmanande körförhållandena på Buffalo-Pittsburgh Highway, och passerar ofta genom isolerad obygdsterräng.
Om du inte är van vid att köra på landsvägar, håll huvudet kallt: branta lutningar, smala körfält och skarpa kurvor dominerar.
Skyltade hastighetsbegränsningar är märkbart lägre än i tidigare och efterföljande avsnitt - vanligtvis 35-40 mph (56-64 km/h) - och strikt lydnad mot dem är ännu viktigare än annars.
Märkligt nog är dock mobiltelefontjänsten mycket starkare här än längs många andra sträckor av rutten, t.ex. Pennsylvania Wilds.
Tyska bakverk är ganska goda, och i Bayern är de ganska rika och varierade, liknande dem i deras södra granne, Österrike.
Fruktbakelser är vanliga, med äpplen som kokas till bakverk året runt, och körsbär och plommon som dyker upp under sommaren.
Många tyska bakverk innehåller också mandel, hasselnötter och andra trädnötter. Populära kakor passar ofta särskilt bra till en kopp starkt kaffe.
Om du vill ha några små men mustiga bakverk kan du prova det som beroende på region kallas Berliner, Pfannkuchen eller Krapfen.
En curry är en maträtt baserad på örter och kryddor, tillsammans med antingen kött eller grönsaker.
En curry kan vara antingen "torr" eller "våt" beroende på mängden vätska.
I inlandsregionerna i norra Indien och Pakistan används yoghurt ofta i curryrätter; I södra Indien och vissa andra kustregioner på subkontinenten används kokosmjölk ofta.
Med 17 000 öar att välja mellan är indonesisk mat ett paraplybegrepp som täcker ett stort utbud av regionala kök som finns över hela landet.
Men om termen används utan ytterligare bestämningar tenderar den att betyda den mat som ursprungligen kommer från de centrala och östra delarna av huvudön Java.
Det javanesiska köket, som nu är allmänt tillgängligt i hela skärgården, har en rad enkelt kryddade rätter, där de dominerande smaksättningarna som javaneserna föredrar är jordnötter, chili, socker (särskilt javanesiskt kokossocker) och olika aromatiska kryddor.
Stigbyglar är stöd för ryttarens fötter som hänger ner på vardera sidan av sadeln.
De ger större stabilitet för ryttaren men kan ha säkerhetsproblem på grund av risken för att en ryttares fötter fastnar i dem.
Om en ryttare kastas av en häst men har en fot som fastnat i stigbygeln kan de dras om hästen springer iväg. För att minimera denna risk kan ett antal säkerhetsåtgärder vidtas.
För det första bär de flesta ryttare ridstövlar med häl och en slät, ganska smal sula.
Därefter har vissa sadlar, särskilt engelska sadlar, säkerhetsstänger som gör att ett stigläder kan falla av sadeln om det dras bakåt av en fallande ryttare.
Cochamó Valley - Chiles främsta klättringsdestination, känd som Sydamerikas Yosemite, med en mängd olika granitväggar och klippor.
Topparna inkluderar hisnande vyer från topparna. Klättrare från alla delar av världen etablerar ständigt nya rutter bland dess oändliga potential av väggar.
Utförsåkningssporter, som inkluderar skidåkning och snowboard, är populära sporter som innebär att man glider nerför snötäckt terräng med skidor eller en snowboard fäst vid fötterna.
Skidåkning är en stor reseaktivitet med många entusiaster, ibland kända som "ski bums", som planerar hela semestrar kring skidåkning på en viss plats.
Idén om skidåkning är mycket gammal - grottmålningar som föreställer skidåkare går tillbaka så långt som 5000 f.Kr.!
Utförsåkning som sport går tillbaka till åtminstone 1600-talet, och 1861 öppnades den första fritidsskidklubben av norrmän i Australien.
Backpacking på skidor: Denna aktivitet kallas också backcountry ski, ski touring eller ski hiking.
Det är relaterat till men involverar vanligtvis inte alpina skidturer eller bergsklättring, de senare görs i brant terräng och kräver mycket styvare skidor och pjäxor.
Tänk på skidrutten som en liknande vandringsled.
Under bra förhållanden kommer du att kunna tillryggalägga något längre sträckor än att gå – men det är mycket sällan du kommer att få längdskidåkningens hastigheter utan en tung ryggsäck i preparerade spår.
Europa är en kontinent som är relativt liten men med många självständiga länder. Under normala omständigheter skulle resor genom flera länder innebära att man måste gå igenom visumansökningar och passkontroll flera gånger.
Schengenområdet fungerar dock lite som ett land i detta avseende.
Så länge du håller dig i denna zon kan du i allmänhet korsa gränserna utan att gå igenom passkontrollerna igen.
På samma sätt, genom att ha ett Schengenvisum, behöver du inte ansöka om visum till vart och ett av Schengenmedlemsländerna separat, vilket sparar tid, pengar och pappersarbete.
Det finns ingen universell definition för vilka tillverkade föremål som är antikviteter. Vissa skatteverk definierar varor som är äldre än 100 år som antikviteter.
Definitionen har geografiska variationer, där åldersgränsen kan vara kortare på platser som Nordamerika än i Europa.
Hantverksprodukter kan definieras som antikviteter, även om de är yngre än liknande massproducerade varor.
Renskötseln är en viktig näring bland samerna och kulturen kring näringen är viktig även för många med andra yrken.
Inte heller traditionellt har alla samer sysslat med storskalig renskötsel, utan livnärt sig på fiske, jakt och liknande, och har renar mest som dragdjur.
Idag arbetar många samer inom moderna yrken. Turismen är en viktig inkomstkälla i det samiska området Sápmi.
Även om ordet "zigenare" används flitigt, särskilt bland icke-romer, anses det ofta stötande på grund av dess associationer till negativa stereotyper och felaktiga uppfattningar om romer.
Om landet du ska besöka blir föremål för en reseavrådan kan din resesjukförsäkring eller din avbeställningsförsäkring påverkas.
Du kanske också vill konsultera råd från andra regeringar än din egen, men deras råd är utformade för deras medborgare.
Som ett exempel kan amerikanska medborgare i Mellanöstern ställas inför andra situationer än européer eller araber.
Bulletiner är bara en kort sammanfattning av den politiska situationen i ett land.
De synpunkter som presenteras är ofta summariska, allmänna och alltför förenklade jämfört med den mer detaljerade information som finns tillgänglig på annat håll.
Hårt väder är den generiska termen för alla farliga väderfenomen med potential att orsaka skada, allvarliga sociala störningar eller förlust av människoliv.
Oväder kan förekomma var som helst i världen, och det finns olika typer av det, som kan bero på geografi, topografi och atmosfäriska förhållanden.
Kraftiga vindar, hagel, kraftig nederbörd och skogsbränder är former och effekter av hårt väder, liksom åskväder, tornados, vattenpip och cykloner.
Regionala och säsongsbetonade ovädersfenomen inkluderar snöstormar, snöstormar, isstormar och sandstormar.
Resenärer rekommenderas starkt att vara medvetna om eventuella risker för hårt väder som påverkar deras område eftersom de kan påverka alla resplaner.
Den som planerar ett besök i ett land som kan betraktas som en krigszon bör få professionell utbildning.
En sökning på Internet efter "Hostile environment course" kommer förmodligen att ge adressen till ett lokalt företag.
En kurs kommer normalt att täcka alla de frågor som diskuteras här mycket mer i detalj, vanligtvis med praktisk erfarenhet.
En kurs kommer normalt att vara från 2-5 dagar och kommer att innebära rollspel, mycket första hjälpen och ibland vapenträning.
Böcker och tidskrifter som handlar om överlevnad i vildmarken är vanliga, men publikationer som handlar om krigszoner är få.
Resenärer som planerar könsbyteskirurgi utomlands måste se till att de har med sig giltiga dokument för återresan.
Regeringarnas vilja att utfärda pass med kön som inte anges (X) eller dokument som uppdaterats för att matcha ett önskat namn och kön varierar.
Utländska regeringars beredvillighet att respektera dessa dokument varierar lika mycket.
Genomsökningar vid säkerhetskontroller har också blivit mycket mer påträngande efter den 11 september 2001.
Transpersoner som inte opererar ska inte förvänta sig att passera genom skannrar med sin integritet och värdighet i behåll.
Ripströmmar är det återkommande flödet från vågor som bryter från stranden, ofta vid ett rev eller liknande.
På grund av undervattenstopologin är returflödet koncentrerat till några djupare sektioner, och en snabb ström till djupt vatten kan bildas där.
De flesta dödsfall inträffar till följd av trötthet när man försöker simma tillbaka mot strömmen, vilket kan vara omöjligt.
Så fort du kommer ut ur strömmen är det inte svårare att simma tillbaka än normalt.
Försök att sikta någonstans där du inte fångas igen eller, beroende på dina färdigheter och om du har blivit upptäckt, kanske du vill vänta på räddning.
Återinträdeschocken kommer tidigare än kulturchocken (det finns mindre av en smekmånadsfas), varar längre och kan vara allvarligare.
Resenärer som hade lätt att anpassa sig till den nya kulturen har ibland särskilt svårt att anpassa sig till sin ursprungskultur.
När du återvänder hem efter att ha bott utomlands har du anpassat dig till den nya kulturen och förlorat några av dina vanor från din hemkultur.
När du åkte utomlands i början var folk förmodligen tålmodiga och förstående, eftersom de visste att resenärer i ett nytt land måste anpassa sig.
Människor kanske inte förväntar sig att tålamod och förståelse också är nödvändigt för resenärer som återvänder hem.
Pyramidens ljud- och ljusshow är en av de mest intressanta sakerna i området för barn.
Du kan se pyramiderna i mörkret och du kan se dem i tystnad innan föreställningen börjar.
Vanligtvis hör du alltid ljudet av turister och försäljare. Berättelsen om ljud och ljus är precis som en sagobok.
Sfinxen är satt som bakgrund och berättare i en lång berättelse.
Scenerna visas på pyramiderna och de olika pyramiderna är upplysta.
Sydshetlandsöarna, som upptäcktes 1819, hävdas av flera nationer och har flest baser, med sexton aktiva 2020.
Skärgården ligger 120 km norr om halvön. Den största är King George Island med bosättningen Villa Las Estrellas.
Andra inkluderar Livingston Island och Deception där den översvämmade kalderan av en fortfarande aktiv vulkan ger en spektakulär naturhamn.
Ellsworth Land är regionen söder om halvön, avgränsad av Bellingshausenhavet.
Bergen på halvön smälter samman med platån och återuppstår sedan för att bilda den 360 km långa kedjan av Ellsworth Mountains, som delas av Minnesotaglaciären.
Den norra delen eller Sentinel Range har Antarktis högsta berg, Vinsonmassivet, som toppar på 4892 m Mount Vinson.
På avlägsna platser, utan mobiltelefontäckning, kan en satellittelefon vara ditt enda alternativ.
En satellittelefon är i allmänhet inte en ersättning för en mobiltelefon, eftersom du måste vara utomhus med fri sikt till satelliten för att ringa ett telefonsamtal.
Tjänsten används ofta av sjöfarten, inklusive fritidsbåtar, samt expeditioner som har behov av fjärrdata och röst.
Din lokala telefonleverantör bör kunna ge mer information om hur du ansluter till den här tjänsten.
Ett allt populärare alternativ för dem som planerar ett sabbatsår är att resa och lära sig.
Detta är särskilt populärt bland dem som lämnar skolan, vilket gör att de kan ta ett sabbatsår före universitetet utan att kompromissa med sin utbildning.
I många fall kan en sabbatsårskurs utomlands faktiskt förbättra dina chanser att komma in på högre utbildning i ditt hemland.
Vanligtvis kommer det att finnas en studieavgift för att anmäla sig till dessa utbildningsprogram.
Finland är en utmärkt båtdestination. "De tusen sjöarnas land" har också tusentals öar, i sjöarna och i kustskärgårdarna.
I skärgårdar och sjöar behöver du inte nödvändigtvis en yacht.
Även om kustskärgårdarna och de största sjöarna verkligen är tillräckligt stora för alla yachter, erbjuder mindre båtar eller till och med en kajak en annan upplevelse.
Båtliv är ett nationellt tidsfördriv i Finland, med en båt till var sjunde eller åttonde person.
Detta matchas av Norge, Sverige och Nya Zeeland, men annars är det ganska unikt (t.ex. i Nederländerna är siffran en till fyrtio).
De flesta av de distinkta Östersjökryssningarna har en längre vistelse i Sankt Petersburg, Ryssland.
Det betyder att du kan besöka den historiska staden i ett par hela dagar medan du återvänder och sover på fartyget på natten.
Om du bara går i land med hjälp av utflykter ombord behöver du inget separat visum (från och med 2009).
Vissa kryssningar har Berlin, Tyskland i broschyrerna. Som du kan se på kartan ovan ligger Berlin inte i närheten av havet och ett besök i staden ingår inte i priset för kryssningen.
Att resa med flyg kan vara en skrämmande upplevelse för människor i alla åldrar och bakgrunder, särskilt om de inte har flugit tidigare eller har upplevt en traumatisk händelse.
Det är inte något att skämmas för: det skiljer sig inte från de personliga rädslor och motpoler mot andra saker som väldigt många människor har.
För vissa kan förståelse för hur flygplan fungerar och vad som händer under en flygning hjälpa till att övervinna en rädsla som bygger på det okända eller på att man inte har kontroll.
Budfirmor får bra betalt för att leverera saker snabbt. Ofta är tiden mycket viktig med affärsdokument, varor eller reservdelar för en brådskande reparation.
På vissa rutter har de större bolagen egna flygplan, men för andra rutter och mindre företag fanns det ett problem.
Om de skickade saker med flygfrakt kan det på vissa rutter ha tagit dagar att komma igenom lossning och tull.
Det enda sättet att få igenom den snabbare var att skicka den som incheckat bagage. Flygbolagens regler tillåter dem inte att skicka bagage utan passagerare, och det är där du kommer in.
Det självklara sättet att flyga i första klass eller business class är att punga ut med en tjock bunt pengar för privilegiet (eller, ännu bättre, få ditt företag att göra det åt dig).
Detta är dock inte billigt: som grova tumregler kan du räkna med att betala upp till fyra gånger det normala ekonomipriset för affärer och elva gånger för första klass!
Generellt sett är det ingen idé att ens leta efter rabatter för affärs- eller förstaklassplatser på direktflyg från A till B.
Flygbolagen vet mycket väl att det finns en viss kärngrupp av flygare som är villiga att betala dyra pengar för privilegiet att komma någonstans snabbt och bekvämt, och ta betalt därefter.
Moldaviens huvudstad är Chisinau. Det lokala språket är rumänska, men ryska används i stor utsträckning.
Moldavien är en multietnisk republik som har drabbats av etniska konflikter.
1994 ledde denna konflikt till skapandet av den självutnämnda republiken Transnistrien i östra Moldavien, som har en egen regering och valuta men som inte erkänns av något av FN:s medlemsländer.
De ekonomiska banden har återupprättats mellan dessa två delar av Moldavien trots att de politiska förhandlingarna har misslyckats.
Den största religionen i Moldavien är ortodoxt kristen.
İzmir är den tredje största staden i Turkiet med en befolkning på cirka 3,7 miljoner, den näst största hamnen efter Istanbul och ett mycket bra transportnav.
En gång i tiden var det den antika staden Smyrna, men nu är det ett modernt, utvecklat och livligt kommersiellt centrum, som ligger runt en enorm bukt och omges av berg.
De breda boulevarderna, byggnaderna med glasfasader och moderna köpcentrum är översållade med traditionella röda tegeltak, 1700-talsmarknaden och gamla moskéer och kyrkor, även om staden har en atmosfär som är mer av medelhavseuropa än det traditionella Turkiet.
Byn Haldarsvík erbjuder utsikt över den närliggande ön Eysturoy och har en ovanlig åttkantig kyrka.
På kyrkogården finns intressanta marmorskulpturer av duvor över några gravar.
Det är värt en halvtimme att strosa runt i den spännande byn.
I norr och inom räckhåll ligger den romantiska och fascinerande staden Sintra och som blev känd för utlänningar efter en glödande berättelse om dess prakt nedtecknad av Lord Byron.
Scotturb Bus 403 går regelbundet till Sintra och stannar vid Cabo da Roca.
I norr kan du också besöka den stora helgedomen Vår Fru av Fatima (helgedomen), en plats för världsberömda Mariauppenbarelser.
Kom ihåg att du i huvudsak besöker en massgravplats, såväl som en plats som har en nästan oberäknelig betydelse för en betydande del av världens befolkning.
Det finns fortfarande många män och kvinnor i livet som överlevde sin tid här, och många fler som hade nära och kära som mördades eller arbetade ihjäl sig där, både judar och icke-judar.
Behandla webbplatsen med all den värdighet, högtidlighet och respekt den förtjänar. Skämta inte om Förintelsen eller nazister.
Förstör inte platsen genom att markera eller repa graffiti i strukturer.
Barcelonas officiella språk är katalanska och spanska. Ungefär hälften föredrar att tala katalanska, en stor majoritet förstår det och i stort sett alla kan spanska.
De flesta skyltar anges dock endast på katalanska eftersom det är fastställt i lag som det första officiella språket.
Men spanska används också i stor utsträckning i kollektivtrafiken och andra anläggningar.
Regelbundna meddelanden i tunnelbanan görs endast på katalanska, men oplanerade störningar meddelas av ett automatiserat system på en mängd olika språk, inklusive spanska, engelska, franska, arabiska och japanska.
Parisarna har ett rykte om sig att vara egocentriska, oförskämda och arroganta.
Även om detta ofta bara är en felaktig stereotyp, är det bästa sättet att komma överens i Paris fortfarande att uppföra sig på bästa sätt och bete sig som någon som är "bien élevé" (väl uppfostrad). Det kommer att göra det betydligt lättare att ta sig fram.
Parisarnas plötsliga yttre kommer snabbt att försvinna om du visar några grundläggande artigheter.
Nationalparken Plitvicesjöarna är kraftigt skogbevuxen, främst med bok, gran och gran, och har en blandning av alpin och medelhavsvegetation.
Den har en anmärkningsvärt stor variation av växtsamhällen på grund av dess varierande mikroklimat, olika jordar och varierande nivåer av höjd.
Området är också hem för en mycket stor variation av djur- och fågelarter.
Sällsynta djur som brunbjörn, varg, örn, uggla, lodjur, vildkatt och tjäder finns där, tillsammans med många vanligare arter
När kvinnor besöker klostren måste de bära kjolar som täcker knäna och ha axlarna täckta.
De flesta av klostren tillhandahåller wraps för kvinnor som kommer oförberedda, men om du tar med dig din egen, särskilt en med ljusa färger, får du ett leende från munken eller nunnan vid ingången.
På samma sätt måste män bära byxor som täcker knäna.
Även detta kan lånas från lagret vid entrén men de kläderna tvättas inte efter varje användare så du kanske inte känner dig bekväm med att bära dessa kjolar. En storlek passar alla för män!
Det mallorkinska köket, liksom det i liknande områden i Medelhavet, är baserat på bröd, grönsaker och kött (särskilt fläskkött) och använder olivolja genomgående.
En enkel populär middag, särskilt under sommaren, är Pa amb Oli: Bröd med olivolja, tomat och alla tillgängliga kryddor som ost, tonfisk etc.
Alla substantiv, tillsammans med ordet Sie för dig, börjar alltid med stor bokstav, även mitt i en mening.
Detta är ett viktigt sätt att skilja mellan vissa verb och objekt.
Det gör det också lättare att läsa, även om skrivandet är något komplicerat av behovet av att ta reda på om ett verb eller adjektiv används i en substantiviserad form.
Uttalet är relativt enkelt på italienska eftersom de flesta ord uttalas exakt som de skrivs
De viktigaste bokstäverna att se upp för är c och g, eftersom deras uttal varierar beroende på följande vokal.
Se också till att uttala r och rr på olika sätt: caro betyder kär, medan carro betyder vagn.
Persiska har en relativt lätt och mestadels regelbunden grammatik.
Att läsa denna grammatikprimer skulle därför hjälpa dig att lära dig mycket om persisk grammatik och förstå fraser bättre.
Det behöver inte sägas att om du kan ett romanskt språk blir det lättare för dig att lära dig portugisiska.
Men människor som kan lite spanska kan snabbt dra slutsatsen att portugisiskan är tillräckligt nära för att den inte behöver studeras separat.
Förmoderna observatorier är vanligtvis föråldrade idag och finns kvar som museer eller utbildningsplatser.
Eftersom ljusföroreningar under deras storhetstid inte var den typ av problem som det är idag, är de vanligtvis belägna i städer eller på campus, lättare att nå än de som byggdes i modern tid.
De flesta moderna forskningsteleskop är enorma anläggningar i avlägsna områden med gynnsamma atmosfäriska förhållanden.
Att titta på körsbärsblommor, känd som hanami, har varit en del av den japanska kulturen sedan 700-talet.
Konceptet kom från Kina där plommonblommor var den blomma som gällde.
I Japan anordnade kejsaren de första körsbärsblomsfesterna endast för sig själv och andra medlemmar av aristokratin runt det kejserliga hovet.
Växter ser bäst ut när de befinner sig i en naturlig miljö, så motstå frestelsen att ta bort även "bara ett" exemplar.
Om du besöker en formellt arrangerad trädgård kommer du också att bli utkastad utan diskussion om du samlar in "exemplar".
Singapore är i allmänhet en extremt säker plats att vara på och mycket lätt att navigera, och du kan köpa nästan vad som helst efter ankomsten.
Men eftersom du befinner dig i de "höga tropikerna" bara några grader norr om ekvatorn måste du hantera både värme (alltid) och stark sol (när himlen är klar, mer sällan).
Det finns också några bussar som går norrut till Hebron, den traditionella begravningsplatsen för de bibliska patriarkerna Abraham, Isak, Jakob och deras fruar.
Kontrollera att bussen du funderar på att ta går in till Hebron och inte bara till den närliggande judiska bosättningen Kiryat Arba.
Inre vattenvägar kan vara ett bra tema att basera en semester kring.
Till exempel besöka slott i Loiredalen, Rhendalen eller ta en kryssning till intressanta städer vid Donau eller åka båt längs Eriekanalen.
De definierar också rutter för populära vandrings- och cykelleder.
Julen är en av kristendomens viktigaste högtider och firas som Jesu födelsedag.
Många av traditionerna kring högtiden har också anammats av icke-troende i kristna länder och icke-kristna runt om i världen.
Det finns en tradition att tillbringa påsknatten vaken vid någon exponerad punkt för att se soluppgången.
Det finns naturligtvis kristna teologiska förklaringar till denna tradition, men det kan mycket väl vara en förkristen vår- och fruktbarhetsritual.
Mer traditionella kyrkor håller ofta en påskvaka på lördagskvällen under påskhelgen, och församlingarna bryter ofta ut i firande vid tolvslaget, för att fira Kristi uppståndelse.
Alla djur som ursprungligen anlände till öarna kom hit antingen genom att simma, flyga eller flyta.
På grund av det långa avståndet från kontinenten kunde däggdjur inte göra resan, vilket gjorde jättesköldpaddan till det primära betesdjuret på Galapagos.
Sedan människans ankomst till Galapagos har många däggdjur introducerats, bland annat getter, hästar, kor, råttor, katter och hundar.
Om du besöker Arktis eller Antarktis på vintern kommer du att uppleva polarnatten, vilket innebär att solen inte går upp över horisonten.
Detta ger ett bra tillfälle att se norrskenet, eftersom himlen kommer att vara mörk mer eller mindre dygnet runt.
Eftersom områdena är glest befolkade och ljusföroreningar därför ofta inte är ett problem, kommer du också att kunna njuta av stjärnorna.
Den japanska arbetskulturen är mer hierarkisk och formell än vad västerlänningar kanske är vana vid.
Kostymer är vanliga affärskläder och medarbetare kallar varandra vid efternamn eller jobbtitlar.
Harmoni på arbetsplatsen är avgörande, med betoning på gruppinsatser snarare än att berömma individuella prestationer.
Arbetstagare måste ofta få sina överordnades godkännande för alla beslut de fattar, och förväntas lyda sina överordnades instruktioner utan att ifrågasätta.
